# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

##################################################################################
#
#           GLOBALFOUNDRIES
#
##################################################################################
#
# 180MCU Tech LEF File
# based on DRM DM-000013-01 Rev 13
# TFG-Version: 2.1.9
# Date: February 2018
#-------------------------------------------------------
# metal stack option: 5LM_1TM_11K
# Preferred routing directions:
# vertical:   Metal2 Metal4 
# horizontal: Metal1 Metal3 Metal5
#------------------------------------------------------
# This Techfile contains not correct Parasitic Information.
# USE Appropriate parasitic files for Parasitic Extraction.
#------------------------------------------------------

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
    DATABASE MICRONS 2000  ;
    CAPACITANCE PICOFARADS 1 ;
    CURRENT MILLIAMPS 1 ;
    RESISTANCE OHMS 1 ;
END UNITS

SITE GF018hv5v_green_sc9
  SYMMETRY X Y ;
  CLASS core ;
  SIZE 0.56 BY 5.04 ;
END GF018hv5v_green_sc9

PROPERTYDEFINITIONS
  LAYER LEF58_EOLENCLOSURE STRING ;
  LAYER LEF58_TYPE STRING ;
END PROPERTYDEFINITIONS

MANUFACTURINGGRID 0.0050 ;
CLEARANCEMEASURE EUCLIDEAN ;
USEMINSPACING OBS ON ;

LAYER Pwell
    TYPE MASTERSLICE ;
    PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
END Pwell

LAYER Nwell
    TYPE MASTERSLICE ;
    PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
END Nwell

LAYER Poly2
    TYPE MASTERSLICE ;
END Poly2

LAYER CON
    TYPE CUT ;
END CON



LAYER Metal1
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;

    PITCH 0.56 ;
    OFFSET 0.0 ;  

    MINWIDTH 0.230 ;                   # Mn.1  (n=1)
    WIDTH 0.230 ;                      # Mn.1  (n=1)
    SPACING 0.230  ;                   # Mn.2a (n=1)
    SPACING 0.300 RANGE 10.005 999.00 ; # Mn.2b
    AREA 0.1444 ;                      # Mn.3

    THICKNESS 0.54 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNASIDEAREARATIO 400 ;

    DCCURRENTDENSITY AVERAGE 0.67 ;
    ACCURRENTDENSITY AVERAGE 1.00 ;

    CAPACITANCE CPERSQDIST 0.0004 ;
    RESISTANCE RPERSQ 0.090 ;

    MINIMUMDENSITY 30.0 ;
    DENSITYCHECKWINDOW 200.0 200.0 ;
    DENSITYCHECKSTEP 100.0 ;

END Metal1


LAYER Via1
  TYPE CUT ;
  SPACING 0.26 ;
  WIDTH   0.26 ;

  ENCLOSURE BELOW 0.00 0.06 ;
  ENCLOSURE ABOVE 0.01 0.06 ;
  PROPERTY LEF58_EOLENCLOSURE "
  	EOLENCLOSURE 0.34 0.06 ;" ; 

  ARRAYSPACING CUTSPACING 0.36 ARRAYCUTS 4 SPACING 0.36 ; # Vn.2b
  RESISTANCE 4.5 ;

  ACCURRENTDENSITY AVERAGE 0.28 ;
  DCCURRENTDENSITY AVERAGE 0.18 ;
  ANTENNAMODEL OXIDE1 ;
  ANTENNAAREARATIO 20.0 ;
END Via1


LAYER Metal2
    TYPE ROUTING ;
    DIRECTION VERTICAL ;

    PITCH 0.56 ;
    OFFSET 0.0 ;  

    MINWIDTH 0.280 ;
    WIDTH 0.280 ;                        # Mn.1  (n>1)
    SPACING 0.280 ;                      # Mn.2a (n>1)
    SPACING 0.300 RANGE 10.005 999.00 ;  # Mn.2b
    AREA 0.1444 ;                        # Mn.3

    THICKNESS 0.54 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFSIDEAREARATIO 400 ;
    ANTENNAGATEPLUSDIFF 2 ;

    DCCURRENTDENSITY AVERAGE 0.67 ;
    ACCURRENTDENSITY AVERAGE 1.00 ;

    CAPACITANCE CPERSQDIST 0.0003 ;
    RESISTANCE RPERSQ 0.090 ;

    MINIMUMDENSITY 30.0 ;
    DENSITYCHECKWINDOW 200.0 200.0 ;
    DENSITYCHECKSTEP 100.0 ;

END Metal2


LAYER Via2
  TYPE CUT ;
  SPACING 0.26 ;
  WIDTH   0.26 ;

  ENCLOSURE BELOW 0.01 0.06 ;
  ENCLOSURE ABOVE 0.01 0.06 ;

  # a bit conservative for Vn.3/4a without considering the protrusion length of 0.28
  PROPERTY LEF58_EOLENCLOSURE " EOLENCLOSURE 0.34 0.06 ; " ;

  ARRAYSPACING CUTSPACING 0.36 ARRAYCUTS 4 SPACING 0.36 ; # Vn.2b
  RESISTANCE 4.5 ;

  ACCURRENTDENSITY AVERAGE 0.28 ;
  DCCURRENTDENSITY AVERAGE 0.18 ;
  ANTENNAMODEL OXIDE1 ;
  ANTENNAAREARATIO 20.0 ;
END Via2


LAYER Metal3
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;

    PITCH 0.56 ;
    OFFSET 0.0 ;  

    MINWIDTH 0.280 ;
    WIDTH 0.280 ;                        # Mn.1  (n>1)
    SPACING 0.280 ;                      # Mn.2a (n>1)
    SPACING 0.300 RANGE 10.005 999.00 ;  # Mn.2b
    AREA 0.1444 ;                        # Mn.3

    THICKNESS 0.54 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFSIDEAREARATIO 400 ;
    ANTENNAGATEPLUSDIFF 2 ;

    DCCURRENTDENSITY AVERAGE 0.67 ;
    ACCURRENTDENSITY AVERAGE 1.00 ;

    CAPACITANCE CPERSQDIST 0.00028 ;
    RESISTANCE RPERSQ 0.090 ;

    MINIMUMDENSITY 30.0 ;
    DENSITYCHECKWINDOW 200.0 200.0 ;
    DENSITYCHECKSTEP 100.0 ;

END Metal3


LAYER Via3
  TYPE CUT ;
  SPACING 0.26 ;
  WIDTH   0.26 ;

  ENCLOSURE BELOW 0.01 0.06 ;
  ENCLOSURE ABOVE 0.01 0.06 ;

  # a bit conservative for Vn.3/4a without considering the protrusion length of 0.28
  PROPERTY LEF58_EOLENCLOSURE " EOLENCLOSURE 0.34 0.06 ; " ;

  ARRAYSPACING CUTSPACING 0.36 ARRAYCUTS 4 SPACING 0.36 ; # Vn.2b
  RESISTANCE 4.5 ;

  ACCURRENTDENSITY AVERAGE 0.28 ;
  DCCURRENTDENSITY AVERAGE 0.18 ;
  ANTENNAMODEL OXIDE1 ;
  ANTENNAAREARATIO 20.0 ;
END Via3


LAYER Metal4
    TYPE ROUTING ;
    DIRECTION VERTICAL ;

    PITCH 0.56 ;
    OFFSET 0.0 ;  

    MINWIDTH 0.280 ;
    WIDTH 0.280 ;                        # Mn.1  (n>1)
    SPACING 0.280 ;                      # Mn.2a (n>1)
    SPACING 0.300 RANGE 10.005 999.00 ;  # Mn.2b
    AREA 0.1444 ;                        # Mn.3

    THICKNESS 0.54 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFSIDEAREARATIO 400 ;
    ANTENNAGATEPLUSDIFF 2 ;

    DCCURRENTDENSITY AVERAGE 0.67 ;
    ACCURRENTDENSITY AVERAGE 1.00 ;

    CAPACITANCE CPERSQDIST 0.000277 ;
    RESISTANCE RPERSQ 0.090 ;

    MINIMUMDENSITY 30.0 ;
    DENSITYCHECKWINDOW 200.0 200.0 ;
    DENSITYCHECKSTEP 100.0 ;

END Metal4


LAYER Via4
  TYPE CUT ;
  SPACING 0.26 ;
  WIDTH   0.26 ;

  ENCLOSURE BELOW 0.01 0.06 ;
  ENCLOSURE ABOVE 0.01 0.06 ;

  # a bit conservative for Vn.3/4a without considering the protrusion length of 0.28
  PROPERTY LEF58_EOLENCLOSURE " EOLENCLOSURE 0.34 0.06 ; " ;

  ARRAYSPACING CUTSPACING 0.36 ARRAYCUTS 4 SPACING 0.36 ; # Vn.2b
  RESISTANCE 4.5 ;

  ACCURRENTDENSITY AVERAGE 0.28 ;
  DCCURRENTDENSITY AVERAGE 0.18 ;
  ANTENNAMODEL OXIDE1 ;
  ANTENNAAREARATIO 20.0 ;
END Via4



LAYER Metal5
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;

    OFFSET 0.0 ;  


    PITCH 0.9 ;
    MINWIDTH 0.440 ;
    WIDTH   0.440 ;                      # MT.1
    AREA    0.5625 ;                     # MT.4
    SPACING 0.460 ;                      # MT.2a
    SPACING 0.600 RANGE 10.005 999.00 ;  # MT.2b

    DCCURRENTDENSITY AVERAGE 1.5 ;
    ACCURRENTDENSITY AVERAGE 2.2 ;
    RESISTANCE RPERSQ 0.060 ;

    THICKNESS 1.19 ;

    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFSIDEAREARATIO 400 ;
    ANTENNAGATEPLUSDIFF 2 ;

    CAPACITANCE CPERSQDIST 0.0000394 ;

    MINIMUMDENSITY 30.0 ;
    DENSITYCHECKWINDOW 200.0 200.0 ;
    DENSITYCHECKSTEP 100.0 ;

END Metal5



LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

LAYER PR_bndry
    TYPE MASTERSLICE ;
END PR_bndry


#------------------------------------------------------------
#  Via1 VIA SECTION 
#------------------------------------------------------------
 VIA Via1_HH  DEFAULT
 LAYER Via1 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal1 ;
 RECT -0.190 -0.130 0.190 0.130 ;
 LAYER Metal2 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 RESISTANCE 4.500 ;
 END Via1_HH 
 
 VIA Via1_HV  DEFAULT
 LAYER Via1 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal1 ;
 RECT -0.190 -0.130 0.190 0.130 ;
 LAYER Metal2 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 RESISTANCE 4.500 ;
 END Via1_HV 
 
 VIA Via1_VH  DEFAULT
 LAYER Via1 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal1 ;
 RECT -0.130 -0.190 0.130 0.190 ;
 LAYER Metal2 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 RESISTANCE 4.500 ;
 END Via1_VH 
 
 VIA Via1_VV  DEFAULT
 LAYER Via1 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal1 ;
 RECT -0.130 -0.190 0.130 0.190 ;
 LAYER Metal2 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 RESISTANCE 4.500 ;
 END Via1_VV 
 
 VIA Via1_2CUT_H
 LAYER Via1 ;
 RECT -0.390 -0.130 -0.130 0.130 ;
 RECT 0.130 -0.130 0.390 0.130 ;
 LAYER Metal1 ;
 RECT -0.450 -0.130 0.450 0.130 ;
 LAYER Metal2 ;
 RECT -0.400 -0.190 0.400 0.190 ;
 END Via1_2CUT_H
 
 VIA Via1_2CUT_V
 LAYER Via1 ;
 RECT -0.130 -0.390 0.130 -0.130 ;
 RECT -0.130 0.130 0.130 0.390 ;
 LAYER Metal1 ;
 RECT -0.190 -0.390 0.190 0.390 ;
 LAYER Metal2 ;
 RECT -0.140 -0.450 0.140 0.450 ;
 END Via1_2CUT_V
 
 VIA Via1_2X2_0_60_10_60_H_H  DEFAULT
 LAYER Via1 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal1 ;
 RECT -0.450 -0.390 0.450 0.390 ;
 LAYER Metal2 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 END Via1_2X2_0_60_10_60_H_H 
 
 VIA Via1_2X2_0_60_10_60_H_V  DEFAULT
 LAYER Via1 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal1 ;
 RECT -0.450 -0.390 0.450 0.390 ;
 LAYER Metal2 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 END Via1_2X2_0_60_10_60_H_V 
 
 VIA Via1_2X2_0_60_10_60_V_H  DEFAULT
 LAYER Via1 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal1 ;
 RECT -0.390 -0.450 0.390 0.450 ;
 LAYER Metal2 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 END Via1_2X2_0_60_10_60_V_H 
 
 VIA Via1_2X2_0_60_10_60_V_V  DEFAULT
 LAYER Via1 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal1 ;
 RECT -0.390 -0.450 0.390 0.450 ;
 LAYER Metal2 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 END Via1_2X2_0_60_10_60_V_V 
 
VIARULE Via1_GEN_HH GENERATE
  LAYER Metal1 ;
    ENCLOSURE 0.060 0.000 ;
  LAYER Metal2 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER Via1 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via1_GEN_HH

VIARULE Via1_GEN_HV GENERATE
  LAYER Metal1 ;
    ENCLOSURE 0.060 0.000 ;
  LAYER Metal2 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER Via1 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via1_GEN_HV

VIARULE Via1_GEN_VH GENERATE
  LAYER Metal1 ;
    ENCLOSURE 0.000 0.060 ;
  LAYER Metal2 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER Via1 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via1_GEN_VH

VIARULE Via1_GEN_VV GENERATE
  LAYER Metal1 ;
    ENCLOSURE 0.000 0.060 ;
  LAYER Metal2 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER Via1 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via1_GEN_VV

 VIA Via1_4X4H_HH_DEFAULT  DEFAULT
 LAYER Via1 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal1 ;
 RECT -1.120 -1.060 1.120 1.060 ;
 LAYER Metal2 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 END Via1_4X4H_HH_DEFAULT 
 
 VIA Via1_4X4H_HV_DEFAULT  DEFAULT
 LAYER Via1 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal1 ;
 RECT -1.120 -1.060 1.120 1.060 ;
 LAYER Metal2 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 END Via1_4X4H_HV_DEFAULT 
 
 VIA Via1_4X4H_VH_DEFAULT  DEFAULT
 LAYER Via1 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal1 ;
 RECT -1.060 -1.120 1.060 1.120 ;
 LAYER Metal2 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 END Via1_4X4H_VH_DEFAULT 
 
 VIA Via1_4X4H_VV_DEFAULT  DEFAULT
 LAYER Via1 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal1 ;
 RECT -1.060 -1.120 1.060 1.120 ;
 LAYER Metal2 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 END Via1_4X4H_VV_DEFAULT 
 
#------------------------------------------------------------
#  Via2 VIA SECTION 
#------------------------------------------------------------
 VIA Via2_HH  DEFAULT
 LAYER Via2 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal2 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 LAYER Metal3 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 RESISTANCE 4.500 ;
 END Via2_HH 
 
 VIA Via2_HV  DEFAULT
 LAYER Via2 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal2 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 LAYER Metal3 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 RESISTANCE 4.500 ;
 END Via2_HV 
 
 VIA Via2_VH  DEFAULT
 LAYER Via2 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal2 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 LAYER Metal3 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 RESISTANCE 4.500 ;
 END Via2_VH 
 
 VIA Via2_VV  DEFAULT
 LAYER Via2 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal2 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 LAYER Metal3 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 RESISTANCE 4.500 ;
 END Via2_VV 
 
 VIA Via2_2CUT_H
 LAYER Via2 ;
 RECT -0.390 -0.130 -0.130 0.130 ;
 RECT 0.130 -0.130 0.390 0.130 ;
 LAYER Metal2 ;
 RECT -0.390 -0.190 0.390 0.190 ;
 LAYER Metal3 ;
 RECT -0.450 -0.140 0.450 0.140 ;
 END Via2_2CUT_H
 
 VIA Via2_2CUT_V
 LAYER Via2 ;
 RECT -0.130 -0.390 0.130 -0.130 ;
 RECT -0.130 0.130 0.130 0.390 ;
 LAYER Metal2 ;
 RECT -0.130 -0.450 0.130 0.450 ;
 LAYER Metal3 ;
 RECT -0.190 -0.400 0.190 0.400 ;
 END Via2_2CUT_V
 
 VIA Via2_2X2_0_60_10_60_H_H  DEFAULT
 LAYER Via2 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal2 ;
 RECT -0.450 -0.390 0.450 0.390 ;
 LAYER Metal3 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 END Via2_2X2_0_60_10_60_H_H 
 
 VIA Via2_2X2_0_60_10_60_H_V  DEFAULT
 LAYER Via2 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal2 ;
 RECT -0.450 -0.390 0.450 0.390 ;
 LAYER Metal3 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 END Via2_2X2_0_60_10_60_H_V 
 
 VIA Via2_2X2_0_60_10_60_V_H  DEFAULT
 LAYER Via2 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal2 ;
 RECT -0.390 -0.450 0.390 0.450 ;
 LAYER Metal3 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 END Via2_2X2_0_60_10_60_V_H 
 
 VIA Via2_2X2_0_60_10_60_V_V  DEFAULT
 LAYER Via2 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal2 ;
 RECT -0.390 -0.450 0.390 0.450 ;
 LAYER Metal3 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 END Via2_2X2_0_60_10_60_V_V 
 
VIARULE Via2_GEN_HH GENERATE
  LAYER Metal2 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER Metal3 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER Via2 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via2_GEN_HH

VIARULE Via2_GEN_HV GENERATE
  LAYER Metal2 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER Metal3 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER Via2 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via2_GEN_HV

VIARULE Via2_GEN_VH GENERATE
  LAYER Metal2 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER Metal3 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER Via2 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via2_GEN_VH

VIARULE Via2_GEN_VV GENERATE
  LAYER Metal2 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER Metal3 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER Via2 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via2_GEN_VV

 VIA Via2_4X4H_HH_DEFAULT  DEFAULT
 LAYER Via2 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal2 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 LAYER Metal3 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 END Via2_4X4H_HH_DEFAULT 
 
 VIA Via2_4X4H_HV_DEFAULT  DEFAULT
 LAYER Via2 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal2 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 LAYER Metal3 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 END Via2_4X4H_HV_DEFAULT 
 
 VIA Via2_4X4H_VH_DEFAULT  DEFAULT
 LAYER Via2 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal2 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 LAYER Metal3 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 END Via2_4X4H_VH_DEFAULT 
 
 VIA Via2_4X4H_VV_DEFAULT  DEFAULT
 LAYER Via2 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal2 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 LAYER Metal3 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 END Via2_4X4H_VV_DEFAULT 
 
#------------------------------------------------------------
#  Via3 VIA SECTION 
#------------------------------------------------------------
 VIA Via3_HH  DEFAULT
 LAYER Via3 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal3 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 LAYER Metal4 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 RESISTANCE 4.500 ;
 END Via3_HH 
 
 VIA Via3_HV  DEFAULT
 LAYER Via3 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal3 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 LAYER Metal4 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 RESISTANCE 4.500 ;
 END Via3_HV 
 
 VIA Via3_VH  DEFAULT
 LAYER Via3 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal3 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 LAYER Metal4 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 RESISTANCE 4.500 ;
 END Via3_VH 
 
 VIA Via3_VV  DEFAULT
 LAYER Via3 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal3 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 LAYER Metal4 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 RESISTANCE 4.500 ;
 END Via3_VV 
 
 VIA Via3_2CUT_H
 LAYER Via3 ;
 RECT -0.390 -0.130 -0.130 0.130 ;
 RECT 0.130 -0.130 0.390 0.130 ;
 LAYER Metal3 ;
 RECT -0.450 -0.130 0.450 0.130 ;
 LAYER Metal4 ;
 RECT -0.400 -0.190 0.400 0.190 ;
 END Via3_2CUT_H
 
 VIA Via3_2CUT_V
 LAYER Via3 ;
 RECT -0.130 -0.390 0.130 -0.130 ;
 RECT -0.130 0.130 0.130 0.390 ;
 LAYER Metal3 ;
 RECT -0.190 -0.390 0.190 0.390 ;
 LAYER Metal4 ;
 RECT -0.140 -0.450 0.140 0.450 ;
 END Via3_2CUT_V
 
 VIA Via3_2X2_0_60_10_60_H_H  DEFAULT
 LAYER Via3 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal3 ;
 RECT -0.450 -0.390 0.450 0.390 ;
 LAYER Metal4 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 END Via3_2X2_0_60_10_60_H_H 
 
 VIA Via3_2X2_0_60_10_60_H_V  DEFAULT
 LAYER Via3 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal3 ;
 RECT -0.450 -0.390 0.450 0.390 ;
 LAYER Metal4 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 END Via3_2X2_0_60_10_60_H_V 
 
 VIA Via3_2X2_0_60_10_60_V_H  DEFAULT
 LAYER Via3 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal3 ;
 RECT -0.390 -0.450 0.390 0.450 ;
 LAYER Metal4 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 END Via3_2X2_0_60_10_60_V_H 
 
 VIA Via3_2X2_0_60_10_60_V_V  DEFAULT
 LAYER Via3 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal3 ;
 RECT -0.390 -0.450 0.390 0.450 ;
 LAYER Metal4 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 END Via3_2X2_0_60_10_60_V_V 
 
VIARULE Via3_GEN_HH GENERATE
  LAYER Metal3 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER Metal4 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER Via3 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via3_GEN_HH

VIARULE Via3_GEN_HV GENERATE
  LAYER Metal3 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER Metal4 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER Via3 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via3_GEN_HV

VIARULE Via3_GEN_VH GENERATE
  LAYER Metal3 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER Metal4 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER Via3 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via3_GEN_VH

VIARULE Via3_GEN_VV GENERATE
  LAYER Metal3 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER Metal4 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER Via3 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via3_GEN_VV

 VIA Via3_4X4H_HH_DEFAULT  DEFAULT
 LAYER Via3 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal3 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 LAYER Metal4 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 END Via3_4X4H_HH_DEFAULT 
 
 VIA Via3_4X4H_HV_DEFAULT  DEFAULT
 LAYER Via3 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal3 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 LAYER Metal4 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 END Via3_4X4H_HV_DEFAULT 
 
 VIA Via3_4X4H_VH_DEFAULT  DEFAULT
 LAYER Via3 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal3 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 LAYER Metal4 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 END Via3_4X4H_VH_DEFAULT 
 
 VIA Via3_4X4H_VV_DEFAULT  DEFAULT
 LAYER Via3 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal3 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 LAYER Metal4 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 END Via3_4X4H_VV_DEFAULT 
 
#------------------------------------------------------------
#  Via4 VIA SECTION 
#------------------------------------------------------------
 VIA Via4_HH  DEFAULT
 LAYER Via4 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal4 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 LAYER Metal5 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 RESISTANCE 4.500 ;
 END Via4_HH 
 
 VIA Via4_HV  DEFAULT
 LAYER Via4 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal4 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 LAYER Metal5 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 RESISTANCE 4.500 ;
 END Via4_HV 
 
 VIA Via4_VH  DEFAULT
 LAYER Via4 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal4 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 LAYER Metal5 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 RESISTANCE 4.500 ;
 END Via4_VH 
 
 VIA Via4_VV  DEFAULT
 LAYER Via4 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal4 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 LAYER Metal5 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 RESISTANCE 4.500 ;
 END Via4_VV 
 
 VIA Via4_2CUT_H
 LAYER Via4 ;
 RECT -0.390 -0.130 -0.130 0.130 ;
 RECT 0.130 -0.130 0.390 0.130 ;
 LAYER Metal4 ;
 RECT -0.400 -0.190 0.400 0.190 ;
 LAYER Metal5 ;
 RECT -0.450 -0.140 0.450 0.140 ;
 END Via4_2CUT_H
 
 VIA Via4_2CUT_V
 LAYER Via4 ;
 RECT -0.130 -0.390 0.130 -0.130 ;
 RECT -0.130 0.130 0.130 0.390 ;
 LAYER Metal4 ;
 RECT -0.140 -0.450 0.140 0.450 ;
 LAYER Metal5 ;
 RECT -0.190 -0.400 0.190 0.400 ;
 END Via4_2CUT_V
 
 VIA Via4_2X2_10_60_10_60_H_H  DEFAULT
 LAYER Via4 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal4 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 LAYER Metal5 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 END Via4_2X2_10_60_10_60_H_H 
 
 VIA Via4_2X2_10_60_10_60_H_V  DEFAULT
 LAYER Via4 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal4 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 LAYER Metal5 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 END Via4_2X2_10_60_10_60_H_V 
 
 VIA Via4_2X2_10_60_10_60_V_H  DEFAULT
 LAYER Via4 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal4 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 LAYER Metal5 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 END Via4_2X2_10_60_10_60_V_H 
 
 VIA Via4_2X2_10_60_10_60_V_V  DEFAULT
 LAYER Via4 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal4 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 LAYER Metal5 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 END Via4_2X2_10_60_10_60_V_V 
 
VIARULE Via4_GEN_HH GENERATE
  LAYER Metal4 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER Metal5 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER Via4 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via4_GEN_HH

VIARULE Via4_GEN_HV GENERATE
  LAYER Metal4 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER Metal5 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER Via4 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via4_GEN_HV

VIARULE Via4_GEN_VH GENERATE
  LAYER Metal4 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER Metal5 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER Via4 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via4_GEN_VH

VIARULE Via4_GEN_VV GENERATE
  LAYER Metal4 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER Metal5 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER Via4 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via4_GEN_VV

 VIA Via4_4X4H_HH_DEFAULT  DEFAULT
 LAYER Via4 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal4 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 LAYER Metal5 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 END Via4_4X4H_HH_DEFAULT 
 
 VIA Via4_4X4H_HV_DEFAULT  DEFAULT
 LAYER Via4 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal4 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 LAYER Metal5 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 END Via4_4X4H_HV_DEFAULT 
 
 VIA Via4_4X4H_VH_DEFAULT  DEFAULT
 LAYER Via4 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal4 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 LAYER Metal5 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 END Via4_4X4H_VH_DEFAULT 
 
 VIA Via4_4X4H_VV_DEFAULT  DEFAULT
 LAYER Via4 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal4 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 LAYER Metal5 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 END Via4_4X4H_VV_DEFAULT 
 


MACRO gf180mcu_fd_sc_mcu9t5v0__addf_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addf_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.800 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.265 2.330 3.455 2.710 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.525 2.265 13.850 2.710 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.547000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.890 2.115 12.550 2.345 ;
        RECT 11.910 1.770 12.170 2.115 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.830 2.890 16.475 3.685 ;
        RECT 16.145 0.845 16.475 2.890 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.324400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 0.845 0.575 3.830 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 16.800 5.490 ;
        RECT 1.365 3.875 1.595 4.590 ;
        RECT 6.625 3.610 6.855 4.590 ;
        RECT 8.665 3.140 8.895 4.590 ;
        RECT 10.705 3.505 10.935 4.590 ;
        RECT 15.125 3.875 15.355 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 17.230 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 17.230 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.305 ;
        RECT 6.625 0.450 6.855 1.425 ;
        RECT 8.865 0.450 9.095 1.425 ;
        RECT 10.705 0.450 10.935 1.425 ;
        RECT 15.125 0.450 15.355 1.165 ;
        RECT 0.000 -0.450 16.800 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 4.385 3.170 4.615 3.790 ;
        RECT 1.805 2.940 4.615 3.170 ;
        RECT 5.605 3.265 5.835 3.845 ;
        RECT 9.685 3.265 9.915 3.845 ;
        RECT 11.725 3.265 11.955 3.845 ;
        RECT 5.605 3.035 7.930 3.265 ;
        RECT 9.685 3.035 11.955 3.265 ;
        RECT 12.845 3.170 13.075 3.685 ;
        RECT 12.845 2.940 14.310 3.170 ;
        RECT 1.805 2.060 2.035 2.940 ;
        RECT 12.845 2.805 13.075 2.940 ;
        RECT 5.010 2.575 13.075 2.805 ;
        RECT 0.870 1.885 2.035 2.060 ;
        RECT 14.080 2.115 14.310 2.940 ;
        RECT 14.080 2.005 15.795 2.115 ;
        RECT 0.870 1.655 4.615 1.885 ;
        RECT 4.385 1.315 4.615 1.655 ;
        RECT 5.505 1.655 7.975 1.885 ;
        RECT 5.505 1.315 5.735 1.655 ;
        RECT 7.745 1.315 7.975 1.655 ;
        RECT 9.585 1.655 11.680 1.885 ;
        RECT 9.585 1.315 9.815 1.655 ;
        RECT 11.450 1.540 11.680 1.655 ;
        RECT 12.945 1.775 15.795 2.005 ;
        RECT 11.450 1.310 12.110 1.540 ;
        RECT 12.945 1.315 13.175 1.775 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addf_1
MACRO gf180mcu_fd_sc_mcu9t5v0__addf_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addf_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.700000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.425 2.330 4.605 2.710 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.700000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.710 2.150 16.110 2.710 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.525000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.050 1.920 13.850 2.150 ;
        RECT 13.590 1.770 13.850 1.920 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.622400 ;
    PORT
      LAYER Metal1 ;
        RECT 17.165 2.710 17.395 3.685 ;
        RECT 17.165 0.845 17.770 2.710 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.622400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 0.845 1.855 3.830 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 19.040 5.490 ;
        RECT 0.605 3.845 0.835 4.590 ;
        RECT 2.645 3.845 2.875 4.590 ;
        RECT 7.785 3.905 8.015 4.590 ;
        RECT 10.025 3.435 10.255 4.590 ;
        RECT 11.765 3.435 11.995 4.590 ;
        RECT 15.965 3.905 16.195 4.590 ;
        RECT 18.185 3.845 18.415 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 19.470 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 19.470 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.285 0.450 0.515 1.165 ;
        RECT 2.525 0.450 2.755 1.165 ;
        RECT 7.785 0.450 8.015 1.215 ;
        RECT 10.025 0.450 10.255 1.215 ;
        RECT 11.865 0.450 12.095 1.215 ;
        RECT 16.265 0.450 16.495 1.195 ;
        RECT 18.505 0.450 18.735 1.165 ;
        RECT 0.000 -0.450 19.040 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 5.545 3.170 5.775 3.685 ;
        RECT 2.965 2.940 5.775 3.170 ;
        RECT 8.805 3.160 9.035 3.740 ;
        RECT 2.965 2.115 3.195 2.940 ;
        RECT 5.545 2.875 5.775 2.940 ;
        RECT 6.710 2.930 9.035 3.160 ;
        RECT 10.745 3.160 10.975 3.740 ;
        RECT 12.885 3.160 13.115 3.740 ;
        RECT 10.745 2.930 13.115 3.160 ;
        RECT 14.105 2.985 16.935 3.215 ;
        RECT 14.105 2.700 14.335 2.985 ;
        RECT 6.070 2.470 14.335 2.700 ;
        RECT 2.085 1.775 3.195 2.115 ;
        RECT 2.965 1.600 3.195 1.775 ;
        RECT 2.965 1.370 5.830 1.600 ;
        RECT 6.665 1.445 9.135 1.675 ;
        RECT 6.665 1.315 6.895 1.445 ;
        RECT 8.905 1.315 9.135 1.445 ;
        RECT 10.745 1.445 13.215 1.675 ;
        RECT 16.705 1.655 16.935 2.985 ;
        RECT 10.745 1.315 10.975 1.445 ;
        RECT 12.985 1.315 13.215 1.445 ;
        RECT 14.050 1.425 16.935 1.655 ;
        RECT 14.050 1.370 14.390 1.425 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addf_2
MACRO gf180mcu_fd_sc_mcu9t5v0__addf_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addf_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.700000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.705 1.860 6.785 2.710 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.700000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.965 2.330 18.530 2.710 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.525000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.330 1.920 15.990 2.150 ;
        RECT 11.910 1.770 12.170 1.920 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.635 3.105 19.865 3.685 ;
        RECT 21.875 3.105 22.105 3.685 ;
        RECT 19.635 2.875 22.105 3.105 ;
        RECT 20.725 1.655 21.185 2.875 ;
        RECT 19.685 1.425 22.155 1.655 ;
        RECT 19.685 0.845 19.915 1.425 ;
        RECT 21.925 0.845 22.155 1.425 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.815850 ;
    PORT
      LAYER Metal1 ;
        RECT 1.445 3.105 1.675 3.685 ;
        RECT 3.785 3.105 4.015 3.685 ;
        RECT 1.445 2.875 4.015 3.105 ;
        RECT 2.380 1.655 2.840 2.875 ;
        RECT 1.445 1.425 3.915 1.655 ;
        RECT 1.445 0.845 1.675 1.425 ;
        RECT 3.685 0.845 3.915 1.425 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 23.520 5.490 ;
        RECT 0.325 3.875 0.555 4.590 ;
        RECT 2.555 3.875 2.785 4.590 ;
        RECT 4.905 3.875 5.135 4.590 ;
        RECT 10.065 3.905 10.295 4.590 ;
        RECT 12.205 3.435 12.435 4.590 ;
        RECT 14.145 3.435 14.375 4.590 ;
        RECT 18.465 3.875 18.695 4.590 ;
        RECT 20.750 3.875 20.980 4.590 ;
        RECT 22.945 3.875 23.175 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 23.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 23.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.325 0.450 0.555 1.165 ;
        RECT 2.565 0.450 2.795 1.165 ;
        RECT 4.805 0.450 5.035 1.165 ;
        RECT 10.065 0.450 10.295 1.215 ;
        RECT 12.305 0.450 12.535 1.215 ;
        RECT 14.145 0.450 14.375 1.215 ;
        RECT 18.565 0.450 18.795 1.165 ;
        RECT 20.805 0.450 21.035 1.165 ;
        RECT 23.045 0.450 23.275 1.165 ;
        RECT 0.000 -0.450 23.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 7.825 3.170 8.055 3.685 ;
        RECT 5.245 2.940 8.055 3.170 ;
        RECT 4.310 2.060 4.595 2.585 ;
        RECT 5.245 2.060 5.475 2.940 ;
        RECT 7.825 2.875 8.055 2.940 ;
        RECT 9.045 3.160 9.275 3.740 ;
        RECT 13.125 3.160 13.355 3.740 ;
        RECT 15.165 3.160 15.395 3.740 ;
        RECT 16.285 3.170 16.515 3.750 ;
        RECT 9.045 2.930 11.370 3.160 ;
        RECT 13.125 2.930 15.395 3.160 ;
        RECT 15.625 2.940 19.235 3.170 ;
        RECT 15.625 2.700 15.855 2.940 ;
        RECT 8.450 2.470 15.855 2.700 ;
        RECT 4.310 1.830 5.475 2.060 ;
        RECT 19.005 2.005 19.235 2.940 ;
        RECT 5.245 1.545 5.475 1.830 ;
        RECT 16.385 1.775 19.235 2.005 ;
        RECT 5.245 1.315 8.110 1.545 ;
        RECT 8.945 1.445 11.415 1.675 ;
        RECT 8.945 1.315 9.175 1.445 ;
        RECT 11.185 1.315 11.415 1.445 ;
        RECT 13.025 1.445 15.495 1.675 ;
        RECT 13.025 1.315 13.255 1.445 ;
        RECT 15.265 1.315 15.495 1.445 ;
        RECT 16.385 1.315 16.615 1.775 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addf_4
MACRO gf180mcu_fd_sc_mcu9t5v0__addh_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addh_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.285 2.950 6.075 3.270 ;
        RECT 2.285 2.215 2.515 2.950 ;
        RECT 5.845 2.215 6.075 2.950 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 2.270 5.195 2.650 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 0.845 0.575 4.360 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.845 1.590 9.175 4.360 ;
        RECT 8.550 1.210 9.175 1.590 ;
        RECT 8.945 0.845 9.175 1.210 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 9.520 5.490 ;
        RECT 1.365 3.550 1.595 4.590 ;
        RECT 3.645 3.960 3.875 4.590 ;
        RECT 4.385 3.960 4.615 4.590 ;
        RECT 7.645 3.550 7.875 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.350 ;
        RECT 7.645 0.450 7.875 1.355 ;
        RECT 0.000 -0.450 9.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.625 3.730 2.855 4.360 ;
        RECT 6.570 3.960 7.415 4.190 ;
        RECT 1.825 3.500 6.955 3.730 ;
        RECT 1.825 2.555 2.055 3.500 ;
        RECT 0.925 2.215 2.055 2.555 ;
        RECT 6.725 2.500 6.955 3.500 ;
        RECT 7.185 3.320 7.415 3.960 ;
        RECT 7.185 3.090 7.810 3.320 ;
        RECT 7.580 2.555 7.810 3.090 ;
        RECT 6.725 2.270 7.350 2.500 ;
        RECT 1.825 1.300 2.055 2.215 ;
        RECT 7.580 2.215 8.495 2.555 ;
        RECT 7.580 1.985 7.810 2.215 ;
        RECT 5.405 1.755 7.810 1.985 ;
        RECT 1.825 1.070 3.850 1.300 ;
        RECT 4.285 0.910 4.515 1.355 ;
        RECT 5.405 1.140 5.635 1.755 ;
        RECT 6.525 0.910 6.755 1.355 ;
        RECT 4.285 0.680 6.755 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addh_1
MACRO gf180mcu_fd_sc_mcu9t5v0__addh_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addh_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.760 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.610 2.940 6.010 3.170 ;
        RECT 3.610 2.500 3.840 2.940 ;
        RECT 3.030 2.270 3.840 2.500 ;
        RECT 5.750 2.500 6.010 2.940 ;
        RECT 5.750 2.270 7.160 2.500 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.070 2.150 4.330 2.710 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 0.770 1.615 4.355 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.729500 ;
    PORT
      LAYER Metal1 ;
        RECT 9.985 1.590 10.215 4.355 ;
        RECT 9.985 0.770 10.490 1.590 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 11.760 5.490 ;
        RECT 0.315 3.875 0.545 4.590 ;
        RECT 2.455 3.875 2.685 4.590 ;
        RECT 4.545 3.875 4.775 4.590 ;
        RECT 5.365 3.875 5.595 4.590 ;
        RECT 8.865 3.875 9.095 4.590 ;
        RECT 11.055 3.875 11.285 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 12.190 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.190 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.265 0.450 0.495 1.580 ;
        RECT 2.505 0.450 2.735 1.580 ;
        RECT 8.865 0.450 9.095 1.580 ;
        RECT 11.105 0.450 11.335 1.580 ;
        RECT 0.000 -0.450 11.760 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.525 3.630 3.755 4.325 ;
        RECT 7.505 3.875 8.635 4.215 ;
        RECT 2.570 3.400 8.175 3.630 ;
        RECT 2.570 2.665 2.800 3.400 ;
        RECT 2.015 2.385 2.800 2.665 ;
        RECT 2.015 1.855 2.245 2.385 ;
        RECT 7.945 2.040 8.175 3.400 ;
        RECT 4.545 1.810 8.175 2.040 ;
        RECT 8.405 2.645 8.635 3.875 ;
        RECT 8.405 2.270 9.635 2.645 ;
        RECT 4.545 0.770 4.775 1.810 ;
        RECT 5.265 0.910 5.495 1.580 ;
        RECT 8.405 1.570 8.635 2.270 ;
        RECT 9.400 1.835 9.635 2.270 ;
        RECT 6.385 1.340 8.635 1.570 ;
        RECT 6.385 1.140 6.615 1.340 ;
        RECT 7.505 0.910 7.735 1.110 ;
        RECT 5.265 0.680 7.735 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addh_2
MACRO gf180mcu_fd_sc_mcu9t5v0__addh_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addh_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.300000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 2.630 8.080 2.860 ;
        RECT 1.100 2.215 1.330 2.630 ;
        RECT 3.930 2.285 6.450 2.630 ;
        RECT 7.850 2.500 8.080 2.630 ;
        RECT 7.850 2.270 9.860 2.500 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.300000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.770 2.055 3.050 2.400 ;
        RECT 6.680 2.170 7.620 2.400 ;
        RECT 6.680 2.055 6.910 2.170 ;
        RECT 1.770 1.825 6.910 2.055 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.550500 ;
    PORT
      LAYER Metal1 ;
        RECT 12.470 2.985 15.100 3.215 ;
        RECT 12.470 1.595 12.805 2.985 ;
        RECT 12.470 1.365 15.150 1.595 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.660300 ;
    PORT
      LAYER Metal1 ;
        RECT 16.950 3.320 17.235 4.360 ;
        RECT 19.205 3.320 19.435 4.360 ;
        RECT 16.950 2.960 19.435 3.320 ;
        RECT 19.075 1.790 19.435 2.960 ;
        RECT 16.950 1.430 19.575 1.790 ;
        RECT 16.950 0.695 17.335 1.430 ;
        RECT 19.345 0.695 19.575 1.430 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 21.280 5.490 ;
        RECT 0.295 3.550 0.525 4.590 ;
        RECT 2.335 3.550 2.565 4.590 ;
        RECT 4.425 3.550 4.655 4.590 ;
        RECT 7.915 4.010 8.145 4.590 ;
        RECT 11.275 4.010 11.505 4.590 ;
        RECT 13.695 4.010 13.925 4.590 ;
        RECT 15.885 3.550 16.115 4.590 ;
        RECT 18.125 3.550 18.355 4.590 ;
        RECT 20.335 3.550 20.565 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 21.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.200 ;
        RECT 4.425 0.450 4.655 1.595 ;
        RECT 11.505 0.675 11.735 1.125 ;
        RECT 15.985 0.675 16.215 1.200 ;
        RECT 11.505 0.450 16.215 0.675 ;
        RECT 18.225 0.450 18.455 1.200 ;
        RECT 20.465 0.450 20.695 1.200 ;
        RECT 0.000 -0.450 21.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.315 3.320 1.545 4.360 ;
        RECT 3.405 3.320 3.635 4.360 ;
        RECT 5.725 3.780 5.955 4.360 ;
        RECT 10.155 3.780 10.385 4.360 ;
        RECT 5.725 3.550 15.610 3.780 ;
        RECT 0.640 3.090 10.320 3.320 ;
        RECT 0.640 1.595 0.870 3.090 ;
        RECT 10.090 2.500 10.320 3.090 ;
        RECT 15.380 2.555 15.610 3.550 ;
        RECT 10.090 2.270 12.230 2.500 ;
        RECT 15.380 2.215 18.590 2.555 ;
        RECT 0.640 1.365 2.615 1.595 ;
        RECT 2.385 0.695 2.615 1.365 ;
        RECT 6.790 1.355 12.195 1.585 ;
        RECT 11.965 1.135 12.195 1.355 ;
        RECT 15.380 1.135 15.610 2.215 ;
        RECT 5.670 0.845 10.490 1.075 ;
        RECT 11.965 0.905 15.610 1.135 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addh_4
MACRO gf180mcu_fd_sc_mcu9t5v0__and2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.806000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.710 0.970 2.960 ;
        RECT 0.115 2.150 0.970 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.806000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.710 2.060 2.960 ;
        RECT 1.830 2.150 2.715 2.710 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 0.845 3.855 3.685 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 4.480 5.490 ;
        RECT 0.245 4.345 0.475 4.590 ;
        RECT 2.285 4.345 2.515 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.505 0.450 2.735 1.165 ;
        RECT 0.000 -0.450 4.480 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.210 4.115 1.550 4.170 ;
        RECT 1.210 3.885 3.175 4.115 ;
        RECT 2.945 1.625 3.175 3.885 ;
        RECT 0.190 1.395 3.175 1.625 ;
        RECT 0.190 1.370 0.530 1.395 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and2_1
MACRO gf180mcu_fd_sc_mcu9t5v0__and2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.612000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.330 0.970 2.715 ;
        RECT 0.710 1.905 0.970 2.330 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.612000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 2.330 2.090 2.710 ;
        RECT 1.830 1.900 2.090 2.330 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.420 0.845 3.770 3.685 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.040 5.490 ;
        RECT 0.260 3.685 0.490 4.590 ;
        RECT 2.520 3.875 2.750 4.590 ;
        RECT 4.560 3.875 4.790 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 5.470 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 5.470 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.300 0.450 2.530 1.165 ;
        RECT 4.540 0.450 4.770 1.165 ;
        RECT 0.000 -0.450 5.040 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.280 3.170 1.510 3.750 ;
        RECT 1.280 2.940 2.970 3.170 ;
        RECT 2.740 1.655 2.970 2.940 ;
        RECT 0.260 1.425 2.970 1.655 ;
        RECT 0.260 0.845 0.490 1.425 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and2_2
MACRO gf180mcu_fd_sc_mcu9t5v0__and2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.224000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.205 1.210 2.090 2.060 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.224000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.355 2.290 4.030 2.715 ;
        RECT 0.355 1.770 0.970 2.290 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.445 2.790 8.085 3.685 ;
        RECT 7.485 1.600 8.085 2.790 ;
        RECT 5.390 0.900 8.085 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 9.520 5.490 ;
        RECT 0.245 3.875 0.475 4.590 ;
        RECT 2.285 3.875 2.515 4.590 ;
        RECT 4.325 3.875 4.555 4.590 ;
        RECT 6.545 4.230 6.775 4.590 ;
        RECT 8.585 4.225 8.815 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.165 ;
        RECT 4.325 0.450 4.555 1.165 ;
        RECT 6.510 0.450 6.850 0.640 ;
        RECT 8.805 0.450 9.035 1.165 ;
        RECT 0.000 -0.450 9.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.265 3.180 1.495 3.875 ;
        RECT 3.305 3.180 3.535 3.875 ;
        RECT 1.265 2.950 4.995 3.180 ;
        RECT 4.765 2.315 4.995 2.950 ;
        RECT 4.765 1.975 6.465 2.315 ;
        RECT 4.765 1.655 4.995 1.975 ;
        RECT 2.320 1.425 4.995 1.655 ;
        RECT 2.320 0.845 2.550 1.425 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and2_4
MACRO gf180mcu_fd_sc_mcu9t5v0__and3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.761000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 2.740 1.145 3.345 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.761000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.820 2.740 2.725 3.375 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.761000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.565 1.770 2.955 2.150 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.630 0.845 4.995 3.830 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.600 5.490 ;
        RECT 1.265 4.345 1.495 4.590 ;
        RECT 3.645 4.345 3.875 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.645 0.450 3.875 1.350 ;
        RECT 0.000 -0.450 5.600 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 4.115 0.475 4.315 ;
        RECT 2.285 4.115 3.415 4.315 ;
        RECT 0.245 3.885 3.415 4.115 ;
        RECT 3.185 2.115 3.415 3.885 ;
        RECT 3.185 1.775 4.315 2.115 ;
        RECT 0.245 0.980 0.475 1.355 ;
        RECT 3.185 0.980 3.415 1.775 ;
        RECT 0.245 0.750 3.415 0.980 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and3_1
MACRO gf180mcu_fd_sc_mcu9t5v0__and3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.160 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.115 2.150 0.970 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.210 2.150 2.090 2.710 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.390 2.290 3.210 2.710 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.480 0.845 4.890 3.685 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 6.160 5.490 ;
        RECT 1.320 3.875 1.550 4.590 ;
        RECT 3.360 3.875 3.590 4.590 ;
        RECT 5.580 3.875 5.810 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.590 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.590 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.360 0.450 3.590 1.165 ;
        RECT 5.600 0.450 5.830 1.165 ;
        RECT 0.000 -0.450 6.160 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.340 3.530 2.570 4.110 ;
        RECT 0.245 3.300 4.210 3.530 ;
        RECT 3.980 1.920 4.210 3.300 ;
        RECT 0.300 1.690 4.210 1.920 ;
        RECT 0.300 0.845 0.530 1.690 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and3_2
MACRO gf180mcu_fd_sc_mcu9t5v0__and3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.200 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.245 1.730 3.115 2.150 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.790 2.380 5.000 2.610 ;
        RECT 3.995 1.770 5.000 2.380 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.840 6.020 3.070 ;
        RECT 0.150 2.330 0.995 2.840 ;
        RECT 5.785 2.415 6.020 2.840 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.550 2.925 9.930 3.630 ;
        RECT 9.580 1.600 9.930 2.925 ;
        RECT 7.250 0.895 9.930 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 11.200 5.490 ;
        RECT 0.245 3.505 0.475 4.590 ;
        RECT 2.285 3.975 2.515 4.590 ;
        RECT 4.325 3.975 4.555 4.590 ;
        RECT 6.585 3.875 6.815 4.590 ;
        RECT 8.625 3.875 8.855 4.590 ;
        RECT 10.665 3.875 10.895 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 11.630 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 11.630 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.325 0.450 0.555 0.695 ;
        RECT 6.185 0.450 6.415 1.165 ;
        RECT 8.370 0.450 8.710 0.640 ;
        RECT 10.665 0.450 10.895 1.165 ;
        RECT 0.000 -0.450 11.200 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.265 3.530 1.495 4.110 ;
        RECT 3.305 3.530 3.535 4.110 ;
        RECT 5.345 3.530 5.575 4.110 ;
        RECT 1.265 3.300 6.855 3.530 ;
        RECT 6.625 2.310 6.855 3.300 ;
        RECT 6.625 1.970 9.260 2.310 ;
        RECT 6.625 1.625 6.855 1.970 ;
        RECT 5.500 1.520 6.855 1.625 ;
        RECT 3.305 1.395 6.855 1.520 ;
        RECT 3.305 1.290 5.755 1.395 ;
        RECT 3.305 0.710 3.535 1.290 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and3_4
MACRO gf180mcu_fd_sc_mcu9t5v0__and4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.160 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.716000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.115 2.165 0.975 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.716000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.230 1.210 2.090 2.115 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.716000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.320 1.210 3.210 2.115 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.716000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.830 2.330 4.500 2.710 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.190 2.890 6.045 3.685 ;
        RECT 5.585 0.845 6.045 2.890 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 6.160 5.490 ;
        RECT 0.305 3.155 0.535 4.590 ;
        RECT 2.345 3.155 2.575 4.590 ;
        RECT 4.565 4.345 4.795 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.590 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.590 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 4.565 0.450 4.795 1.350 ;
        RECT 0.000 -0.450 6.160 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.325 2.925 1.555 3.215 ;
        RECT 3.365 2.985 4.960 3.215 ;
        RECT 3.365 2.925 3.595 2.985 ;
        RECT 1.325 2.695 3.595 2.925 ;
        RECT 4.730 2.115 4.960 2.985 ;
        RECT 4.730 2.005 5.235 2.115 ;
        RECT 3.440 1.775 5.235 2.005 ;
        RECT 0.305 0.980 0.535 1.355 ;
        RECT 3.440 0.980 3.670 1.775 ;
        RECT 0.305 0.750 3.670 0.980 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and4_1
MACRO gf180mcu_fd_sc_mcu9t5v0__and4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.115 2.150 0.970 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.200 2.150 2.090 2.710 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.320 2.290 3.210 2.710 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.440 2.330 4.330 2.710 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.580 1.725 6.100 3.685 ;
        RECT 5.190 0.845 6.100 1.725 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.280 5.490 ;
        RECT 0.300 3.875 0.530 4.590 ;
        RECT 2.340 4.345 2.570 4.590 ;
        RECT 4.380 3.875 4.610 4.590 ;
        RECT 6.600 3.875 6.830 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 4.380 0.450 4.610 0.695 ;
        RECT 6.620 0.450 6.850 1.165 ;
        RECT 0.000 -0.450 7.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.360 3.765 3.590 4.235 ;
        RECT 1.320 3.645 3.590 3.765 ;
        RECT 1.320 3.415 4.790 3.645 ;
        RECT 4.560 2.720 4.790 3.415 ;
        RECT 4.560 2.380 5.230 2.720 ;
        RECT 4.560 1.600 4.790 2.380 ;
        RECT 0.245 1.370 4.790 1.600 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and4_2
MACRO gf180mcu_fd_sc_mcu9t5v0__and4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.440 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.790 1.770 3.890 2.150 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.825 2.380 4.750 2.610 ;
        RECT 4.520 2.150 4.750 2.380 ;
        RECT 4.520 1.770 6.030 2.150 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.975 1.540 2.145 2.060 ;
        RECT 6.260 1.830 7.105 2.060 ;
        RECT 6.260 1.540 6.490 1.830 ;
        RECT 0.975 1.310 6.490 1.540 ;
        RECT 0.975 1.210 2.090 1.310 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.115 2.840 5.210 3.070 ;
        RECT 0.115 2.330 0.970 2.840 ;
        RECT 4.980 2.700 5.210 2.840 ;
        RECT 4.980 2.470 8.125 2.700 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.540 2.920 12.210 3.640 ;
        RECT 11.770 1.600 12.210 2.920 ;
        RECT 9.485 0.900 12.210 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 13.440 5.490 ;
        RECT 0.260 3.325 0.490 4.590 ;
        RECT 2.300 3.795 2.530 4.590 ;
        RECT 4.340 3.795 4.570 4.590 ;
        RECT 6.380 3.795 6.610 4.590 ;
        RECT 8.420 3.795 8.650 4.590 ;
        RECT 10.640 3.875 10.870 4.590 ;
        RECT 12.680 3.875 12.910 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 13.870 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.870 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.260 0.450 0.490 1.165 ;
        RECT 8.420 0.450 8.650 0.695 ;
        RECT 10.605 0.450 10.945 0.640 ;
        RECT 12.900 0.450 13.130 1.165 ;
        RECT 0.000 -0.450 13.440 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.280 3.530 1.510 4.110 ;
        RECT 3.320 3.530 3.550 4.110 ;
        RECT 5.360 3.530 5.590 4.110 ;
        RECT 1.280 3.430 5.590 3.530 ;
        RECT 7.400 3.430 7.630 4.010 ;
        RECT 1.280 3.300 9.090 3.430 ;
        RECT 5.400 3.200 9.090 3.300 ;
        RECT 8.860 2.315 9.090 3.200 ;
        RECT 8.860 1.975 10.550 2.315 ;
        RECT 8.860 1.260 9.090 1.975 ;
        RECT 6.715 1.080 9.090 1.260 ;
        RECT 4.285 1.030 9.090 1.080 ;
        RECT 4.285 0.850 6.940 1.030 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and4_4
MACRO gf180mcu_fd_sc_mcu9t5v0__antenna
  CLASS core ANTENNACELL ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__antenna ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.120 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNADIFFAREA 0.406800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 1.315 0.475 3.215 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 1.120 5.490 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 1.550 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 1.550 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.450 1.120 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__antenna
MACRO gf180mcu_fd_sc_mcu9t5v0__aoi21_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi21_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.415 2.655 3.270 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.115 2.285 0.970 2.710 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.467000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 1.805 3.780 2.815 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.755600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 2.150 1.495 3.685 ;
        RECT 1.265 1.770 2.515 2.150 ;
        RECT 2.285 0.845 2.515 1.770 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 4.480 5.490 ;
        RECT 3.485 3.875 3.715 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.165 ;
        RECT 3.585 0.450 3.815 1.565 ;
        RECT 0.000 -0.450 4.480 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 4.130 2.515 4.360 ;
        RECT 0.245 3.550 0.475 4.130 ;
        RECT 2.285 3.550 2.515 4.130 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi21_1
MACRO gf180mcu_fd_sc_mcu9t5v0__aoi21_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi21_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 1.755 5.120 2.300 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.410 2.560 6.605 2.790 ;
        RECT 3.410 1.770 3.660 2.560 ;
        RECT 5.690 2.155 6.605 2.560 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.934000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.115 1.665 0.980 2.150 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.287600 ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 3.250 3.700 3.830 ;
        RECT 5.630 3.250 5.860 3.830 ;
        RECT 2.330 3.020 5.860 3.250 ;
        RECT 2.330 1.490 2.715 3.020 ;
        RECT 2.330 1.155 4.920 1.490 ;
        RECT 1.375 0.925 4.920 1.155 ;
        RECT 3.010 0.680 4.920 0.925 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.280 5.490 ;
        RECT 1.330 4.345 1.560 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.310 0.450 0.540 1.165 ;
        RECT 2.550 0.450 2.780 0.695 ;
        RECT 6.650 0.450 6.880 1.165 ;
        RECT 0.000 -0.450 7.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.310 3.765 0.540 4.360 ;
        RECT 2.445 4.060 6.880 4.290 ;
        RECT 2.445 3.765 2.680 4.060 ;
        RECT 0.310 3.480 2.680 3.765 ;
        RECT 4.610 3.480 4.840 4.060 ;
        RECT 6.650 3.480 6.880 4.060 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi21_2
MACRO gf180mcu_fd_sc_mcu9t5v0__aoi21_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi21_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.440 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.615 2.135 2.845 ;
        RECT 0.710 1.570 0.970 2.615 ;
        RECT 1.905 2.420 2.135 2.615 ;
        RECT 5.665 1.570 5.895 2.110 ;
        RECT 0.710 1.325 5.895 1.570 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.430 2.475 8.310 2.710 ;
        RECT 1.200 2.190 1.430 2.385 ;
        RECT 3.430 2.190 4.365 2.475 ;
        RECT 1.200 1.960 4.365 2.190 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.868000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.630 2.330 12.735 2.750 ;
        RECT 12.470 2.150 12.730 2.330 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.136000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.410 3.305 1.695 3.835 ;
        RECT 3.505 3.305 3.735 3.835 ;
        RECT 5.545 3.305 5.775 3.885 ;
        RECT 7.585 3.305 7.815 3.885 ;
        RECT 1.410 3.245 7.815 3.305 ;
        RECT 1.410 3.075 8.830 3.245 ;
        RECT 7.580 3.015 8.830 3.075 ;
        RECT 8.550 2.020 8.830 3.015 ;
        RECT 8.550 2.000 12.075 2.020 ;
        RECT 6.345 1.790 12.075 2.000 ;
        RECT 6.345 1.770 9.835 1.790 ;
        RECT 6.345 1.095 6.575 1.770 ;
        RECT 2.370 0.865 6.575 1.095 ;
        RECT 9.605 0.840 9.835 1.770 ;
        RECT 11.845 0.840 12.075 1.790 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 13.440 5.490 ;
        RECT 9.850 3.935 10.190 4.590 ;
        RECT 11.890 3.935 12.230 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 13.870 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.870 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.465 0.450 0.695 0.690 ;
        RECT 4.330 0.450 4.670 0.635 ;
        RECT 8.305 0.450 8.535 1.085 ;
        RECT 10.725 0.450 10.955 1.560 ;
        RECT 12.965 0.450 13.195 1.560 ;
        RECT 0.000 -0.450 13.440 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.445 4.115 8.880 4.345 ;
        RECT 0.445 3.535 0.675 4.115 ;
        RECT 2.485 3.535 2.715 4.115 ;
        RECT 4.525 3.535 4.755 4.115 ;
        RECT 6.565 3.535 6.795 4.115 ;
        RECT 8.550 3.705 8.880 4.115 ;
        RECT 10.870 3.705 11.210 4.230 ;
        RECT 12.910 3.705 13.250 4.230 ;
        RECT 8.550 3.475 13.250 3.705 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi21_4
MACRO gf180mcu_fd_sc_mcu9t5v0__aoi22_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi22_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.930 1.210 3.830 2.115 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.950 2.330 4.915 2.710 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.250 1.210 2.090 2.115 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.130 2.175 0.980 2.710 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.365 3.355 3.600 3.830 ;
        RECT 2.350 2.855 3.600 3.355 ;
        RECT 2.350 0.845 2.580 2.855 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.040 5.490 ;
        RECT 1.330 3.875 1.560 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 5.470 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 5.470 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.310 0.450 0.540 1.165 ;
        RECT 4.390 0.450 4.620 1.165 ;
        RECT 0.000 -0.450 5.040 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.310 3.645 0.540 4.360 ;
        RECT 1.820 4.060 4.620 4.290 ;
        RECT 1.820 3.645 2.050 4.060 ;
        RECT 0.310 3.410 2.050 3.645 ;
        RECT 4.390 3.480 4.620 4.060 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi22_1
MACRO gf180mcu_fd_sc_mcu9t5v0__aoi22_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi22_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.960 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 1.720 7.210 2.315 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.950 2.560 8.270 2.790 ;
        RECT 4.950 1.830 5.510 2.560 ;
        RECT 7.860 2.180 8.270 2.560 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.650 1.630 2.090 2.060 ;
        RECT 1.220 1.210 2.090 1.630 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.690 2.290 4.030 2.520 ;
        RECT 0.690 1.770 0.970 2.290 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.322200 ;
    PORT
      LAYER Metal1 ;
        RECT 4.345 3.250 5.575 3.830 ;
        RECT 7.385 3.250 7.615 3.830 ;
        RECT 4.345 3.020 7.615 3.250 ;
        RECT 4.345 1.490 4.720 3.020 ;
        RECT 2.320 1.105 2.550 1.490 ;
        RECT 4.340 1.105 4.720 1.490 ;
        RECT 6.365 1.105 6.595 1.490 ;
        RECT 2.320 0.875 6.595 1.105 ;
        RECT 2.320 0.680 2.550 0.875 ;
        RECT 6.365 0.680 6.595 0.875 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 8.960 5.490 ;
        RECT 1.265 3.875 1.495 4.590 ;
        RECT 3.305 3.875 3.535 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.390 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.390 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.165 ;
        RECT 4.270 0.450 4.610 0.640 ;
        RECT 8.405 0.450 8.635 1.165 ;
        RECT 0.000 -0.450 8.960 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.645 0.475 4.225 ;
        RECT 2.285 3.645 2.515 4.225 ;
        RECT 3.795 4.060 8.635 4.290 ;
        RECT 3.795 3.645 4.025 4.060 ;
        RECT 0.245 3.415 4.025 3.645 ;
        RECT 6.365 3.480 6.595 4.060 ;
        RECT 8.405 3.480 8.635 4.060 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi22_2
MACRO gf180mcu_fd_sc_mcu9t5v0__aoi22_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi22_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.360 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.440 2.710 14.415 2.860 ;
        RECT 11.210 2.630 14.415 2.710 ;
        RECT 11.210 2.270 11.660 2.630 ;
        RECT 14.185 2.215 14.415 2.630 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.325 2.000 9.555 2.555 ;
        RECT 12.470 2.000 13.415 2.400 ;
        RECT 9.325 1.770 13.415 2.000 ;
        RECT 13.185 0.910 13.415 1.770 ;
        RECT 16.125 0.910 16.355 2.555 ;
        RECT 13.185 0.680 16.355 0.910 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.810 2.785 4.435 3.015 ;
        RECT 2.810 2.270 3.210 2.785 ;
        RECT 4.205 2.500 4.435 2.785 ;
        RECT 4.205 2.270 6.070 2.500 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.000 0.915 2.555 ;
        RECT 3.745 2.000 3.975 2.555 ;
        RECT 7.485 2.215 7.955 2.555 ;
        RECT 7.485 2.000 7.715 2.215 ;
        RECT 0.150 1.770 7.715 2.000 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.552000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.865 3.310 9.895 3.900 ;
        RECT 11.705 3.320 11.935 3.900 ;
        RECT 13.745 3.320 13.975 3.900 ;
        RECT 15.270 3.320 16.015 3.900 ;
        RECT 11.195 3.315 16.015 3.320 ;
        RECT 10.965 3.310 16.015 3.315 ;
        RECT 8.865 3.090 16.015 3.310 ;
        RECT 8.865 3.080 11.245 3.090 ;
        RECT 8.865 1.985 9.095 3.080 ;
        RECT 7.945 1.755 9.095 1.985 ;
        RECT 7.945 1.540 8.175 1.755 ;
        RECT 2.285 1.310 8.175 1.540 ;
        RECT 8.865 1.540 9.095 1.755 ;
        RECT 2.285 0.730 2.515 1.310 ;
        RECT 6.365 0.730 6.595 1.310 ;
        RECT 8.865 0.730 10.915 1.540 ;
        RECT 14.765 1.140 14.995 3.090 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.360 5.490 ;
        RECT 1.265 3.245 1.495 4.590 ;
        RECT 3.305 3.705 3.535 4.590 ;
        RECT 5.345 3.705 5.575 4.590 ;
        RECT 7.385 3.705 7.615 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 17.790 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 17.790 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.540 ;
        RECT 4.325 0.450 4.555 1.070 ;
        RECT 8.405 0.450 8.635 1.525 ;
        RECT 12.725 0.450 12.955 1.540 ;
        RECT 16.805 0.450 17.035 1.540 ;
        RECT 0.000 -0.450 17.360 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 8.405 4.130 17.035 4.360 ;
        RECT 0.245 3.015 0.475 4.055 ;
        RECT 2.150 3.475 2.515 4.055 ;
        RECT 4.325 3.475 4.555 4.055 ;
        RECT 6.365 3.475 6.595 4.055 ;
        RECT 8.405 3.475 8.635 4.130 ;
        RECT 10.685 3.540 10.915 4.130 ;
        RECT 12.725 3.550 12.955 4.130 ;
        RECT 14.765 3.550 14.995 4.130 ;
        RECT 2.150 3.245 8.635 3.475 ;
        RECT 16.805 3.245 17.035 4.130 ;
        RECT 2.150 3.015 2.380 3.245 ;
        RECT 0.245 2.785 2.380 3.015 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi22_4
MACRO gf180mcu_fd_sc_mcu9t5v0__aoi211_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi211_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.626000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.770 1.210 2.695 2.115 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.626000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.115 1.705 0.970 2.595 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.925 1.615 3.815 2.150 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.045 1.615 4.915 2.150 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.010200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 0.980 1.530 3.830 ;
        RECT 3.050 1.060 4.860 1.290 ;
        RECT 3.050 0.980 3.280 1.060 ;
        RECT 1.270 0.750 3.280 0.980 ;
        RECT 4.630 0.920 4.860 1.060 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.600 5.490 ;
        RECT 4.530 3.875 4.760 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 0.450 0.480 1.300 ;
        RECT 3.510 0.450 3.740 0.830 ;
        RECT 0.000 -0.450 5.600 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.250 4.130 2.520 4.360 ;
        RECT 0.250 3.550 0.480 4.130 ;
        RECT 2.290 3.550 2.520 4.130 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi211_1
MACRO gf180mcu_fd_sc_mcu9t5v0__aoi211_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi211_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.765 1.770 2.955 2.215 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 2.445 3.770 2.775 ;
        RECT 0.630 2.305 1.155 2.445 ;
        RECT 3.510 1.770 3.770 2.445 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.560 2.470 8.430 2.700 ;
        RECT 4.560 1.725 5.450 2.470 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 1.770 7.295 2.150 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.341000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.210 3.400 4.330 3.630 ;
        RECT 4.070 1.525 4.330 3.400 ;
        RECT 2.205 1.495 4.330 1.525 ;
        RECT 2.205 1.265 4.960 1.495 ;
        RECT 2.205 0.715 2.435 1.265 ;
        RECT 4.730 1.160 4.960 1.265 ;
        RECT 4.730 0.930 7.935 1.160 ;
        RECT 5.465 0.695 5.695 0.930 ;
        RECT 7.705 0.790 7.935 0.930 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 9.520 5.490 ;
        RECT 6.505 4.345 6.735 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.170 ;
        RECT 4.165 0.450 4.395 0.700 ;
        RECT 6.585 0.450 6.815 0.700 ;
        RECT 8.825 0.450 9.055 0.700 ;
        RECT 0.000 -0.450 9.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.860 8.815 4.090 ;
        RECT 0.245 3.280 0.475 3.860 ;
        RECT 8.585 3.280 8.815 3.860 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi211_2
MACRO gf180mcu_fd_sc_mcu9t5v0__aoi211_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi211_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.160 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 2.150 3.850 2.400 ;
        RECT 5.575 2.170 6.640 2.400 ;
        RECT 3.510 1.985 4.890 2.150 ;
        RECT 5.575 1.985 5.805 2.170 ;
        RECT 3.510 1.755 5.805 1.985 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.545 2.630 8.725 2.860 ;
        RECT 1.545 2.215 1.775 2.630 ;
        RECT 5.115 2.215 5.345 2.630 ;
        RECT 6.870 2.215 8.725 2.630 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.860 2.730 19.450 2.960 ;
        RECT 9.860 2.270 10.200 2.730 ;
        RECT 13.505 2.215 13.735 2.730 ;
        RECT 18.960 2.270 19.450 2.730 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.520 1.985 12.860 2.500 ;
        RECT 14.190 2.270 16.500 2.500 ;
        RECT 14.190 2.150 14.420 2.270 ;
        RECT 13.960 1.985 14.420 2.150 ;
        RECT 12.520 1.755 14.420 1.985 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.682000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.935 3.320 2.165 3.900 ;
        RECT 3.975 3.320 4.205 3.900 ;
        RECT 5.750 3.320 6.245 3.900 ;
        RECT 8.055 3.320 8.285 3.900 ;
        RECT 1.085 3.090 8.285 3.320 ;
        RECT 1.085 1.540 1.315 3.090 ;
        RECT 1.085 1.525 3.040 1.540 ;
        RECT 1.085 1.310 18.670 1.525 ;
        RECT 2.955 1.180 18.670 1.310 ;
        RECT 2.955 0.680 3.185 1.180 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 20.160 5.490 ;
        RECT 11.475 3.650 11.705 4.590 ;
        RECT 16.795 3.650 17.025 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 20.590 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 20.590 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.675 0.450 0.905 1.165 ;
        RECT 4.995 0.450 5.225 0.695 ;
        RECT 9.020 0.450 9.360 0.950 ;
        RECT 11.680 0.450 12.020 0.950 ;
        RECT 14.340 0.450 14.680 0.950 ;
        RECT 17.000 0.450 17.340 0.950 ;
        RECT 19.505 0.450 19.735 1.035 ;
        RECT 0.000 -0.450 20.160 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.915 4.130 9.305 4.360 ;
        RECT 0.915 3.550 1.145 4.130 ;
        RECT 2.955 3.550 3.185 4.130 ;
        RECT 4.995 3.550 5.225 4.130 ;
        RECT 7.035 3.550 7.265 4.130 ;
        RECT 9.075 3.420 9.305 4.130 ;
        RECT 14.135 3.420 14.365 4.360 ;
        RECT 19.455 3.420 19.685 4.360 ;
        RECT 9.075 3.190 19.685 3.420 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi211_4
MACRO gf180mcu_fd_sc_mcu9t5v0__aoi221_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi221_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.160 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.626000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.145 2.865 6.040 3.270 ;
        RECT 5.145 2.415 5.375 2.865 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.626000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 2.165 4.330 2.710 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.626000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.255 1.210 2.090 2.065 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.626000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 2.255 1.015 2.710 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.360 1.670 3.210 2.230 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.184000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.565 1.590 4.795 3.685 ;
        RECT 4.565 1.440 5.915 1.590 ;
        RECT 2.425 1.210 5.915 1.440 ;
        RECT 2.425 1.075 2.655 1.210 ;
        RECT 5.685 0.680 5.915 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 6.160 5.490 ;
        RECT 1.365 3.875 1.595 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.590 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.590 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.285 0.450 0.515 1.300 ;
        RECT 3.725 0.450 3.955 0.980 ;
        RECT 0.000 -0.450 6.160 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.545 4.130 5.815 4.360 ;
        RECT 0.345 3.170 0.575 3.750 ;
        RECT 2.385 3.170 2.615 3.685 ;
        RECT 3.545 3.550 3.775 4.130 ;
        RECT 5.585 3.550 5.815 4.130 ;
        RECT 0.345 2.940 2.615 3.170 ;
        RECT 2.385 2.875 2.615 2.940 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi221_1
MACRO gf180mcu_fd_sc_mcu9t5v0__aoi221_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi221_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.760 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.225 2.470 10.490 2.700 ;
        RECT 10.165 1.210 10.490 2.470 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.240 1.590 8.470 2.115 ;
        RECT 7.300 1.210 8.470 1.590 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.945 1.665 3.845 2.180 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.890 2.440 5.480 2.670 ;
        RECT 4.490 2.205 5.480 2.440 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.715 2.145 1.010 2.785 ;
        RECT 0.715 1.915 2.715 2.145 ;
        RECT 2.485 1.435 2.715 1.915 ;
        RECT 4.630 1.520 6.370 1.750 ;
        RECT 4.630 1.435 4.890 1.520 ;
        RECT 2.485 1.205 4.890 1.435 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.111250 ;
    PORT
      LAYER Metal1 ;
        RECT 7.720 3.250 7.950 3.830 ;
        RECT 9.760 3.250 11.110 3.830 ;
        RECT 6.765 3.020 11.110 3.250 ;
        RECT 0.245 1.455 2.255 1.685 ;
        RECT 0.245 1.315 0.475 1.455 ;
        RECT 2.025 0.975 2.255 1.455 ;
        RECT 6.765 1.290 6.995 3.020 ;
        RECT 5.120 1.060 6.995 1.290 ;
        RECT 5.120 0.975 5.350 1.060 ;
        RECT 2.025 0.745 5.350 0.975 ;
        RECT 6.765 0.920 6.995 1.060 ;
        RECT 10.880 0.845 11.110 3.020 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 11.760 5.490 ;
        RECT 2.330 4.400 2.670 4.590 ;
        RECT 4.390 4.400 4.730 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 12.190 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.190 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 5.580 0.450 5.810 0.830 ;
        RECT 8.920 0.450 9.150 1.300 ;
        RECT 0.000 -0.450 11.760 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 6.665 4.170 11.065 4.290 ;
        RECT 0.345 4.060 11.065 4.170 ;
        RECT 0.345 3.940 6.895 4.060 ;
        RECT 0.345 3.360 0.575 3.940 ;
        RECT 1.365 3.480 5.695 3.710 ;
        RECT 6.665 3.480 6.895 3.940 ;
        RECT 8.740 3.480 8.970 4.060 ;
        RECT 1.365 2.900 1.595 3.480 ;
        RECT 3.405 2.900 3.635 3.480 ;
        RECT 5.465 2.900 5.695 3.480 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi221_2
MACRO gf180mcu_fd_sc_mcu9t5v0__aoi221_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi221_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.400 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.210 2.140 14.550 2.500 ;
        RECT 16.930 2.140 17.270 2.400 ;
        RECT 14.210 1.910 17.270 2.140 ;
        RECT 19.540 2.370 21.450 2.600 ;
        RECT 19.540 1.950 19.770 2.370 ;
        RECT 16.950 1.440 17.270 1.910 ;
        RECT 18.000 1.720 19.770 1.950 ;
        RECT 18.000 1.440 18.230 1.720 ;
        RECT 16.950 1.210 18.230 1.440 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.470 2.630 17.740 2.860 ;
        RECT 16.470 2.600 16.700 2.630 ;
        RECT 16.150 2.370 16.700 2.600 ;
        RECT 17.510 2.500 17.740 2.630 ;
        RECT 17.510 2.270 19.310 2.500 ;
        RECT 17.510 1.770 17.770 2.270 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.700 2.085 1.040 2.600 ;
        RECT 3.695 2.085 3.925 2.400 ;
        RECT 0.700 1.985 3.925 2.085 ;
        RECT 6.195 2.370 8.160 2.600 ;
        RECT 6.195 1.985 6.425 2.370 ;
        RECT 0.700 1.855 6.425 1.985 ;
        RECT 3.510 1.755 6.425 1.855 ;
        RECT 3.510 1.210 3.770 1.755 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 2.630 5.965 2.860 ;
        RECT 1.270 2.315 1.985 2.630 ;
        RECT 5.735 2.215 5.965 2.630 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.110 2.270 9.650 2.710 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 8.064500 ;
    PORT
      LAYER Metal1 ;
        RECT 14.605 3.320 14.835 3.900 ;
        RECT 16.645 3.320 16.875 3.900 ;
        RECT 18.685 3.320 18.915 3.900 ;
        RECT 20.725 3.320 20.955 3.900 ;
        RECT 13.590 3.090 20.955 3.320 ;
        RECT 0.245 1.395 3.280 1.625 ;
        RECT 13.590 1.480 13.850 3.090 ;
        RECT 0.245 0.680 0.475 1.395 ;
        RECT 3.050 0.965 3.280 1.395 ;
        RECT 4.430 1.250 16.720 1.480 ;
        RECT 4.430 0.965 4.660 1.250 ;
        RECT 3.050 0.735 4.660 0.965 ;
        RECT 8.555 0.680 8.785 1.250 ;
        RECT 11.165 0.680 11.395 1.250 ;
        RECT 13.405 0.680 13.635 1.250 ;
        RECT 16.490 0.965 16.720 1.250 ;
        RECT 18.460 1.260 21.975 1.490 ;
        RECT 18.460 0.965 18.690 1.260 ;
        RECT 16.490 0.735 18.690 0.965 ;
        RECT 21.745 0.680 21.975 1.260 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 22.400 5.490 ;
        RECT 0.295 3.090 0.525 4.590 ;
        RECT 2.335 3.550 2.565 4.590 ;
        RECT 4.375 3.550 4.605 4.590 ;
        RECT 6.415 3.550 6.645 4.590 ;
        RECT 8.455 3.550 8.685 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 22.830 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 22.830 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.335 0.450 2.565 1.165 ;
        RECT 6.415 0.450 6.645 1.020 ;
        RECT 10.045 0.450 10.275 1.020 ;
        RECT 12.285 0.450 12.515 1.020 ;
        RECT 15.625 0.450 15.855 1.020 ;
        RECT 19.705 0.450 19.935 1.020 ;
        RECT 0.000 -0.450 22.400 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 9.175 4.130 21.975 4.360 ;
        RECT 1.315 3.320 1.545 3.900 ;
        RECT 3.355 3.320 3.585 3.900 ;
        RECT 5.395 3.320 5.625 3.900 ;
        RECT 7.435 3.320 7.665 3.900 ;
        RECT 9.175 3.550 9.405 4.130 ;
        RECT 10.195 3.320 10.425 3.900 ;
        RECT 11.215 3.535 11.445 4.130 ;
        RECT 1.315 3.305 10.425 3.320 ;
        RECT 12.235 3.305 12.465 3.900 ;
        RECT 13.305 3.545 13.535 4.130 ;
        RECT 15.625 3.550 15.855 4.130 ;
        RECT 17.665 3.550 17.895 4.130 ;
        RECT 19.705 3.550 19.935 4.130 ;
        RECT 1.315 3.090 12.465 3.305 ;
        RECT 21.745 3.090 21.975 4.130 ;
        RECT 10.340 3.075 12.465 3.090 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi221_4
MACRO gf180mcu_fd_sc_mcu9t5v0__aoi222_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi222_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.800 2.415 7.725 3.270 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.145 1.770 6.010 2.150 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.670 1.770 3.830 2.150 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.050 2.255 4.910 2.710 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.220 1.210 2.145 2.060 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.115 2.235 1.070 2.710 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.169200 ;
    PORT
      LAYER Metal1 ;
        RECT 6.220 2.875 6.470 3.215 ;
        RECT 6.240 1.590 6.470 2.875 ;
        RECT 6.240 1.490 7.470 1.590 ;
        RECT 3.160 1.210 7.470 1.490 ;
        RECT 3.160 0.680 3.390 1.210 ;
        RECT 7.240 0.680 7.470 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.840 5.490 ;
        RECT 0.400 3.875 0.630 4.590 ;
        RECT 2.440 3.875 2.670 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 8.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.480 0.450 0.710 1.165 ;
        RECT 5.200 0.450 5.430 0.695 ;
        RECT 0.000 -0.450 7.840 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.160 4.130 7.470 4.360 ;
        RECT 1.365 3.170 1.710 3.700 ;
        RECT 3.160 3.550 3.390 4.130 ;
        RECT 4.125 3.170 4.465 3.810 ;
        RECT 5.200 3.550 7.470 4.130 ;
        RECT 1.365 2.940 4.465 3.170 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi222_1
MACRO gf180mcu_fd_sc_mcu9t5v0__aoi222_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi222_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.000 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.700 2.345 12.960 2.575 ;
        RECT 11.775 1.210 12.960 2.345 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.945 1.210 11.050 2.115 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.605 2.380 8.810 2.610 ;
        RECT 7.605 1.770 8.810 2.380 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.255 1.770 6.770 2.150 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.115 2.645 0.970 3.270 ;
        RECT 0.115 2.415 4.065 2.645 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.825 1.770 2.090 2.150 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.275800 ;
    PORT
      LAYER Metal1 ;
        RECT 10.195 3.105 10.425 3.685 ;
        RECT 12.235 3.105 12.465 3.685 ;
        RECT 9.040 2.875 13.485 3.105 ;
        RECT 9.040 1.490 9.470 2.875 ;
        RECT 0.280 0.925 9.470 1.490 ;
        RECT 0.280 0.680 0.510 0.925 ;
        RECT 4.980 0.680 5.210 0.925 ;
        RECT 9.160 0.845 9.470 0.925 ;
        RECT 13.255 0.845 13.485 2.875 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.000 5.490 ;
        RECT 0.280 3.875 0.510 4.590 ;
        RECT 2.320 3.875 2.550 4.590 ;
        RECT 4.360 3.875 4.590 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.430 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.430 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.320 0.450 2.550 0.695 ;
        RECT 7.120 0.450 7.350 0.695 ;
        RECT 11.215 0.450 11.445 0.695 ;
        RECT 0.000 -0.450 14.000 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 5.080 3.915 13.485 4.145 ;
        RECT 1.300 3.105 1.530 3.685 ;
        RECT 3.340 3.105 3.570 3.685 ;
        RECT 5.080 3.335 5.310 3.915 ;
        RECT 6.100 3.105 6.330 3.685 ;
        RECT 7.120 3.335 7.350 3.915 ;
        RECT 8.140 3.105 8.370 3.685 ;
        RECT 9.160 3.335 9.390 3.915 ;
        RECT 11.215 3.335 11.445 3.915 ;
        RECT 13.255 3.335 13.485 3.915 ;
        RECT 1.300 2.875 8.370 3.105 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi222_2
MACRO gf180mcu_fd_sc_mcu9t5v0__aoi222_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi222_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.320 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 17.865 2.150 18.095 2.555 ;
        RECT 17.865 1.985 19.450 2.150 ;
        RECT 20.785 1.985 21.015 2.400 ;
        RECT 24.865 1.985 25.095 2.555 ;
        RECT 17.865 1.755 25.095 1.985 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 20.135 2.770 22.780 2.860 ;
        RECT 19.750 2.630 23.055 2.770 ;
        RECT 19.750 2.270 20.320 2.630 ;
        RECT 22.595 2.215 23.055 2.630 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.670 1.600 9.930 2.555 ;
        RECT 12.625 1.655 12.855 2.400 ;
        RECT 16.605 1.655 16.835 2.555 ;
        RECT 12.625 1.600 16.835 1.655 ;
        RECT 9.670 1.425 16.835 1.600 ;
        RECT 9.670 1.370 12.775 1.425 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.100 2.770 14.140 2.860 ;
        RECT 12.100 2.630 14.895 2.770 ;
        RECT 12.100 2.500 12.330 2.630 ;
        RECT 13.955 2.540 14.895 2.630 ;
        RECT 11.690 1.830 12.330 2.500 ;
        RECT 14.665 2.215 14.895 2.540 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.825 1.985 1.055 2.555 ;
        RECT 3.745 1.985 3.975 2.555 ;
        RECT 7.825 2.150 8.055 2.555 ;
        RECT 6.310 1.985 8.055 2.150 ;
        RECT 0.825 1.755 8.055 1.985 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.285 2.855 5.710 3.015 ;
        RECT 3.285 2.785 6.015 2.855 ;
        RECT 1.830 2.445 2.090 2.710 ;
        RECT 3.285 2.445 3.515 2.785 ;
        RECT 5.490 2.625 6.015 2.785 ;
        RECT 1.830 2.215 3.515 2.445 ;
        RECT 5.785 2.215 6.015 2.625 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.284400 ;
    PORT
      LAYER Metal1 ;
        RECT 18.305 3.230 18.535 3.900 ;
        RECT 20.345 3.320 20.575 3.900 ;
        RECT 22.385 3.320 22.615 3.900 ;
        RECT 19.740 3.230 23.220 3.320 ;
        RECT 24.425 3.230 24.655 3.900 ;
        RECT 17.665 3.090 24.655 3.230 ;
        RECT 17.665 3.015 19.925 3.090 ;
        RECT 17.285 3.000 19.925 3.015 ;
        RECT 23.035 3.000 24.655 3.090 ;
        RECT 17.285 2.785 17.895 3.000 ;
        RECT 17.285 1.195 17.515 2.785 ;
        RECT 0.190 1.140 8.690 1.195 ;
        RECT 17.285 1.155 25.730 1.195 ;
        RECT 13.405 1.140 25.730 1.155 ;
        RECT 0.190 0.925 25.730 1.140 ;
        RECT 0.190 0.910 13.490 0.925 ;
        RECT 24.730 0.710 25.730 0.925 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 26.320 5.490 ;
        RECT 0.245 3.245 0.475 4.590 ;
        RECT 2.285 3.705 2.515 4.590 ;
        RECT 4.325 3.705 4.555 4.590 ;
        RECT 6.365 3.560 6.595 4.590 ;
        RECT 8.405 3.545 8.635 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 26.750 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 26.750 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.230 0.450 2.570 0.680 ;
        RECT 6.310 0.450 6.650 0.680 ;
        RECT 11.110 0.450 11.450 0.680 ;
        RECT 15.245 0.450 15.475 0.695 ;
        RECT 19.325 0.450 19.555 0.695 ;
        RECT 23.405 0.450 23.635 0.695 ;
        RECT 0.000 -0.450 26.320 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 9.125 4.130 25.675 4.360 ;
        RECT 1.265 3.475 1.495 4.055 ;
        RECT 3.305 3.475 3.535 4.055 ;
        RECT 5.345 3.475 5.575 4.055 ;
        RECT 1.265 3.315 6.150 3.475 ;
        RECT 7.385 3.315 7.615 4.055 ;
        RECT 9.125 3.545 9.355 4.130 ;
        RECT 10.145 3.320 10.375 3.900 ;
        RECT 11.165 3.550 11.395 4.130 ;
        RECT 12.185 3.320 12.415 3.900 ;
        RECT 13.205 3.550 13.435 4.130 ;
        RECT 14.225 3.320 14.510 3.900 ;
        RECT 15.245 3.460 15.475 4.130 ;
        RECT 9.405 3.315 14.510 3.320 ;
        RECT 1.265 3.245 14.510 3.315 ;
        RECT 5.930 3.230 14.510 3.245 ;
        RECT 16.265 3.230 16.495 3.900 ;
        RECT 17.285 3.405 17.515 4.130 ;
        RECT 19.325 3.460 19.555 4.130 ;
        RECT 21.365 3.550 21.595 4.130 ;
        RECT 23.405 3.460 23.635 4.130 ;
        RECT 25.445 3.245 25.675 4.130 ;
        RECT 5.930 3.090 16.495 3.230 ;
        RECT 5.930 3.085 9.455 3.090 ;
        RECT 14.325 3.000 16.495 3.090 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi222_4
MACRO gf180mcu_fd_sc_mcu9t5v0__buf_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.853500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 1.015 2.710 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.390 2.890 2.895 3.775 ;
        RECT 2.665 1.590 2.895 2.890 ;
        RECT 2.390 0.740 2.895 1.590 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 3.360 5.490 ;
        RECT 1.365 3.400 1.595 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 3.790 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 3.790 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.080 ;
        RECT 0.000 -0.450 3.360 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.170 0.575 3.775 ;
        RECT 0.345 2.940 2.160 3.170 ;
        RECT 1.930 2.585 2.160 2.940 ;
        RECT 1.930 1.775 2.215 2.585 ;
        RECT 1.930 1.540 2.160 1.775 ;
        RECT 0.245 1.310 2.160 1.540 ;
        RECT 0.245 0.740 0.475 1.310 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_1
MACRO gf180mcu_fd_sc_mcu9t5v0__buf_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.330 0.970 2.710 ;
        RECT 0.630 2.000 0.970 2.330 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.485 3.015 2.715 4.360 ;
        RECT 2.485 2.730 3.280 3.015 ;
        RECT 2.980 1.590 3.280 2.730 ;
        RECT 2.330 1.210 3.280 1.590 ;
        RECT 2.330 0.710 2.715 1.210 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 4.480 5.490 ;
        RECT 1.265 3.550 1.495 4.590 ;
        RECT 3.505 3.550 3.735 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.165 ;
        RECT 3.605 0.450 3.835 1.520 ;
        RECT 0.000 -0.450 4.480 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.320 0.475 4.360 ;
        RECT 0.245 3.090 1.430 3.320 ;
        RECT 1.200 2.500 1.430 3.090 ;
        RECT 1.200 2.270 2.750 2.500 ;
        RECT 1.200 1.625 1.430 2.270 ;
        RECT 0.245 1.395 1.430 1.625 ;
        RECT 0.245 0.710 0.475 1.395 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_2
MACRO gf180mcu_fd_sc_mcu9t5v0__buf_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.585 0.410 2.710 ;
        RECT 0.150 1.770 0.915 2.585 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.207000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.675 3.105 2.905 4.360 ;
        RECT 4.815 3.105 5.045 3.685 ;
        RECT 2.675 2.875 5.045 3.105 ;
        RECT 3.510 2.000 4.005 2.875 ;
        RECT 2.675 1.770 5.145 2.000 ;
        RECT 2.675 0.730 2.905 1.770 ;
        RECT 4.915 0.730 5.145 1.770 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.600 5.490 ;
        RECT 1.265 3.550 1.495 4.590 ;
        RECT 3.695 3.550 3.925 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.555 0.450 1.785 1.165 ;
        RECT 3.795 0.450 4.025 1.540 ;
        RECT 0.000 -0.450 5.600 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.320 0.475 4.360 ;
        RECT 0.245 3.090 1.375 3.320 ;
        RECT 1.145 2.500 1.375 3.090 ;
        RECT 1.145 2.270 3.220 2.500 ;
        RECT 1.145 1.540 1.375 2.270 ;
        RECT 0.245 1.310 1.375 1.540 ;
        RECT 0.245 0.730 0.475 1.310 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_3
MACRO gf180mcu_fd_sc_mcu9t5v0__buf_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 2.270 1.910 2.650 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.605 3.320 3.835 4.360 ;
        RECT 5.745 3.320 6.075 4.360 ;
        RECT 3.605 3.090 6.075 3.320 ;
        RECT 5.575 1.950 6.075 3.090 ;
        RECT 3.605 1.720 6.075 1.950 ;
        RECT 3.605 0.680 3.865 1.720 ;
        RECT 5.845 0.680 6.075 1.720 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.840 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 8.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 6.965 0.450 7.195 1.490 ;
        RECT 0.000 -0.450 7.840 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 1.365 3.090 2.370 3.320 ;
        RECT 2.140 2.500 2.370 3.090 ;
        RECT 2.140 2.270 4.620 2.500 ;
        RECT 2.140 1.920 2.370 2.270 ;
        RECT 1.365 1.690 2.370 1.920 ;
        RECT 1.365 0.680 1.595 1.690 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_4
MACRO gf180mcu_fd_sc_mcu9t5v0__buf_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 2.215 4.205 2.650 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.284000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.845 3.320 6.075 4.360 ;
        RECT 7.985 3.320 8.215 4.360 ;
        RECT 10.225 3.320 10.455 4.360 ;
        RECT 12.465 3.320 12.695 4.360 ;
        RECT 5.845 2.880 12.695 3.320 ;
        RECT 8.970 2.040 9.470 2.880 ;
        RECT 5.845 1.985 9.470 2.040 ;
        RECT 5.845 1.720 12.795 1.985 ;
        RECT 5.845 0.680 6.075 1.720 ;
        RECT 8.055 0.680 8.315 1.720 ;
        RECT 10.325 0.680 10.555 1.720 ;
        RECT 12.565 0.680 12.795 1.720 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.560 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
        RECT 11.345 3.550 11.575 4.590 ;
        RECT 13.585 3.550 13.815 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 6.965 0.450 7.195 1.490 ;
        RECT 9.205 0.450 9.435 1.165 ;
        RECT 11.445 0.450 11.675 1.490 ;
        RECT 13.685 0.450 13.915 1.490 ;
        RECT 0.000 -0.450 14.560 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 3.205 1.595 4.360 ;
        RECT 3.505 3.205 3.735 4.360 ;
        RECT 1.365 2.975 4.665 3.205 ;
        RECT 4.435 2.650 4.665 2.975 ;
        RECT 4.435 2.270 8.740 2.650 ;
        RECT 4.435 1.985 4.665 2.270 ;
        RECT 9.700 2.215 13.220 2.650 ;
        RECT 1.365 1.755 4.665 1.985 ;
        RECT 1.365 0.680 1.595 1.755 ;
        RECT 3.605 0.680 3.835 1.755 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_8
MACRO gf180mcu_fd_sc_mcu9t5v0__buf_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 10.242000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.130 2.270 5.640 2.650 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 10.926000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.135 3.320 8.365 4.360 ;
        RECT 10.275 3.320 10.505 4.360 ;
        RECT 12.515 3.320 12.745 4.360 ;
        RECT 14.755 3.320 14.985 4.360 ;
        RECT 16.995 3.320 17.225 4.360 ;
        RECT 19.235 3.320 19.465 4.360 ;
        RECT 8.135 2.840 19.465 3.320 ;
        RECT 13.500 2.040 14.000 2.840 ;
        RECT 8.135 1.985 14.000 2.040 ;
        RECT 8.135 1.755 19.565 1.985 ;
        RECT 8.135 0.680 8.365 1.755 ;
        RECT 10.375 0.680 10.605 1.755 ;
        RECT 12.385 0.680 12.845 1.755 ;
        RECT 14.855 0.680 15.085 1.755 ;
        RECT 17.095 0.680 17.325 1.755 ;
        RECT 19.335 0.680 19.565 1.755 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 21.280 5.490 ;
        RECT 0.295 3.550 0.525 4.590 ;
        RECT 2.435 3.550 2.665 4.590 ;
        RECT 4.675 3.550 4.905 4.590 ;
        RECT 6.915 3.550 7.145 4.590 ;
        RECT 9.155 3.875 9.385 4.590 ;
        RECT 11.395 3.550 11.625 4.590 ;
        RECT 13.635 3.550 13.865 4.590 ;
        RECT 15.875 3.550 16.105 4.590 ;
        RECT 18.115 3.550 18.345 4.590 ;
        RECT 20.355 3.550 20.585 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 21.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.295 0.450 0.525 1.490 ;
        RECT 2.535 0.450 2.765 1.490 ;
        RECT 4.775 0.450 5.005 1.490 ;
        RECT 7.015 0.450 7.245 1.490 ;
        RECT 9.255 0.450 9.485 1.490 ;
        RECT 11.495 0.450 11.725 1.490 ;
        RECT 13.735 0.450 13.965 1.490 ;
        RECT 15.975 0.450 16.205 1.490 ;
        RECT 18.215 0.450 18.445 1.490 ;
        RECT 20.455 0.450 20.685 1.490 ;
        RECT 0.000 -0.450 21.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.415 3.320 1.645 4.360 ;
        RECT 3.555 3.320 3.785 4.360 ;
        RECT 5.820 3.320 6.225 4.360 ;
        RECT 1.415 2.880 6.225 3.320 ;
        RECT 5.895 2.500 6.225 2.880 ;
        RECT 5.895 2.270 12.910 2.500 ;
        RECT 5.895 2.040 6.225 2.270 ;
        RECT 14.230 2.215 19.630 2.555 ;
        RECT 1.415 1.720 6.225 2.040 ;
        RECT 1.415 0.680 1.645 1.720 ;
        RECT 3.655 0.680 3.885 1.720 ;
        RECT 5.895 0.680 6.225 1.720 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_12
MACRO gf180mcu_fd_sc_mcu9t5v0__buf_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.000 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 13.655999 ;
    PORT
      LAYER Metal1 ;
        RECT 0.440 2.270 7.830 2.650 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 14.568000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.325 3.320 10.555 4.360 ;
        RECT 12.465 3.320 12.695 4.360 ;
        RECT 14.705 3.320 14.935 4.360 ;
        RECT 16.945 3.320 17.175 4.360 ;
        RECT 19.185 3.320 19.415 4.360 ;
        RECT 21.425 3.320 21.655 4.360 ;
        RECT 23.665 3.320 23.895 4.360 ;
        RECT 25.905 3.320 26.135 4.360 ;
        RECT 10.325 2.960 26.135 3.320 ;
        RECT 17.805 2.040 18.555 2.960 ;
        RECT 10.325 1.985 18.555 2.040 ;
        RECT 10.325 1.720 26.235 1.985 ;
        RECT 10.325 0.680 10.555 1.720 ;
        RECT 12.565 0.680 12.795 1.720 ;
        RECT 14.805 0.680 15.035 1.720 ;
        RECT 17.045 0.680 17.305 1.720 ;
        RECT 19.285 0.680 19.515 1.720 ;
        RECT 21.525 0.680 21.755 1.720 ;
        RECT 23.765 0.680 23.995 1.720 ;
        RECT 26.005 0.680 26.235 1.720 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 28.000 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
        RECT 11.345 3.550 11.575 4.590 ;
        RECT 13.585 3.550 13.815 4.590 ;
        RECT 15.825 3.550 16.055 4.590 ;
        RECT 18.065 3.550 18.295 4.590 ;
        RECT 20.305 3.550 20.535 4.590 ;
        RECT 22.545 3.550 22.775 4.590 ;
        RECT 24.785 3.550 25.015 4.590 ;
        RECT 27.025 3.550 27.255 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 28.430 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 28.430 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 6.965 0.450 7.195 1.490 ;
        RECT 9.205 0.450 9.435 1.490 ;
        RECT 11.445 0.450 11.675 1.490 ;
        RECT 13.685 0.450 13.915 1.490 ;
        RECT 15.925 0.450 16.155 1.490 ;
        RECT 18.165 0.450 18.395 1.490 ;
        RECT 20.405 0.450 20.635 1.490 ;
        RECT 22.645 0.450 22.875 1.490 ;
        RECT 24.885 0.450 25.115 1.490 ;
        RECT 27.125 0.450 27.355 1.490 ;
        RECT 0.000 -0.450 28.000 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 5.745 3.320 5.975 4.360 ;
        RECT 8.060 3.320 8.425 4.360 ;
        RECT 1.365 2.880 8.425 3.320 ;
        RECT 8.060 2.630 8.425 2.880 ;
        RECT 8.060 2.270 16.980 2.630 ;
        RECT 8.060 2.040 8.425 2.270 ;
        RECT 18.785 2.215 26.065 2.555 ;
        RECT 1.365 1.720 8.425 2.040 ;
        RECT 1.365 0.680 1.595 1.720 ;
        RECT 3.605 0.680 3.835 1.720 ;
        RECT 5.845 0.680 6.075 1.720 ;
        RECT 8.085 0.680 8.425 1.720 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_16
MACRO gf180mcu_fd_sc_mcu9t5v0__buf_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_20 ;
  ORIGIN 0.000 0.000 ;
  SIZE 34.720 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 17.070000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 2.215 9.845 2.650 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 18.209999 ;
    PORT
      LAYER Metal1 ;
        RECT 12.565 3.320 12.795 4.360 ;
        RECT 14.705 3.320 14.935 4.360 ;
        RECT 16.945 3.320 17.175 4.360 ;
        RECT 19.185 3.320 19.415 4.360 ;
        RECT 21.425 3.320 21.655 4.360 ;
        RECT 23.665 3.320 23.895 4.360 ;
        RECT 25.905 3.320 26.135 4.360 ;
        RECT 28.145 3.320 28.375 4.360 ;
        RECT 30.385 3.320 30.615 4.360 ;
        RECT 32.625 3.320 32.855 4.360 ;
        RECT 12.565 2.885 32.855 3.320 ;
        RECT 22.285 2.880 32.855 2.885 ;
        RECT 22.285 2.030 23.035 2.880 ;
        RECT 12.565 1.980 23.035 2.030 ;
        RECT 12.565 1.720 32.955 1.980 ;
        RECT 12.565 0.680 12.825 1.720 ;
        RECT 14.805 0.680 15.035 1.720 ;
        RECT 17.045 0.680 17.275 1.720 ;
        RECT 19.285 0.680 19.515 1.720 ;
        RECT 21.525 0.680 21.755 1.720 ;
        RECT 23.765 0.680 23.995 1.720 ;
        RECT 26.005 0.680 26.235 1.720 ;
        RECT 28.245 0.680 28.475 1.720 ;
        RECT 30.485 0.680 30.715 1.720 ;
        RECT 32.725 0.680 32.955 1.720 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 34.720 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
        RECT 11.345 3.875 11.575 4.590 ;
        RECT 13.585 3.550 13.815 4.590 ;
        RECT 15.825 3.550 16.055 4.590 ;
        RECT 18.065 3.550 18.295 4.590 ;
        RECT 20.305 3.550 20.535 4.590 ;
        RECT 22.545 3.550 22.775 4.590 ;
        RECT 24.785 3.550 25.015 4.590 ;
        RECT 27.025 3.550 27.255 4.590 ;
        RECT 29.265 3.550 29.495 4.590 ;
        RECT 31.505 3.550 31.735 4.590 ;
        RECT 33.745 3.550 33.975 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 35.150 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 35.150 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 6.965 0.450 7.195 1.490 ;
        RECT 9.205 0.450 9.435 1.490 ;
        RECT 11.445 0.450 11.675 1.490 ;
        RECT 13.685 0.450 13.915 1.490 ;
        RECT 15.925 0.450 16.155 1.490 ;
        RECT 18.165 0.450 18.395 1.490 ;
        RECT 20.405 0.450 20.635 1.490 ;
        RECT 22.645 0.450 22.875 1.490 ;
        RECT 24.885 0.450 25.115 1.490 ;
        RECT 27.125 0.450 27.355 1.490 ;
        RECT 29.365 0.450 29.595 1.490 ;
        RECT 31.605 0.450 31.835 1.490 ;
        RECT 33.845 0.450 34.075 1.490 ;
        RECT 0.000 -0.450 34.720 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 5.745 3.320 5.975 4.360 ;
        RECT 7.985 3.320 8.215 4.360 ;
        RECT 10.225 3.320 10.555 4.360 ;
        RECT 1.365 2.900 10.555 3.320 ;
        RECT 10.225 2.650 10.555 2.900 ;
        RECT 10.225 2.270 21.100 2.650 ;
        RECT 10.225 1.975 10.555 2.270 ;
        RECT 23.265 2.215 32.425 2.650 ;
        RECT 1.365 1.720 10.555 1.975 ;
        RECT 1.365 0.680 1.595 1.720 ;
        RECT 3.605 0.680 3.835 1.720 ;
        RECT 5.845 0.680 6.075 1.720 ;
        RECT 8.085 0.680 8.315 1.720 ;
        RECT 10.325 0.680 10.555 1.720 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_20
MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.698000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.870 2.330 2.090 2.710 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.849000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.630 1.745 4.990 2.150 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.640 1.650 6.870 3.685 ;
        RECT 6.640 0.840 7.130 1.650 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.280 5.490 ;
        RECT 1.365 3.635 1.595 4.590 ;
        RECT 5.440 3.875 5.670 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.425 ;
        RECT 5.660 0.450 5.890 0.690 ;
        RECT 0.000 -0.450 7.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.060 0.575 4.285 ;
        RECT 2.385 4.055 4.650 4.285 ;
        RECT 2.385 3.475 2.615 4.055 ;
        RECT 2.630 2.815 2.895 3.155 ;
        RECT 2.630 2.060 2.860 2.815 ;
        RECT 3.405 2.060 3.635 3.815 ;
        RECT 0.245 1.830 2.860 2.060 ;
        RECT 3.090 1.830 3.635 2.060 ;
        RECT 4.170 2.700 4.650 4.055 ;
        RECT 4.170 2.470 6.345 2.700 ;
        RECT 0.245 1.315 0.475 1.830 ;
        RECT 2.485 0.950 2.715 1.425 ;
        RECT 3.090 1.115 3.320 1.830 ;
        RECT 4.170 1.600 4.400 2.470 ;
        RECT 3.550 1.370 4.400 1.600 ;
        RECT 5.305 1.115 6.385 2.055 ;
        RECT 3.090 0.950 6.385 1.115 ;
        RECT 2.485 0.920 6.385 0.950 ;
        RECT 2.485 0.720 5.430 0.920 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_1
MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.400 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.880 2.330 2.090 2.715 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.692000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.125 2.285 5.465 2.710 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.622400 ;
    PORT
      LAYER Metal1 ;
        RECT 6.705 0.840 7.130 3.720 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 8.400 5.490 ;
        RECT 1.375 3.845 1.605 4.590 ;
        RECT 5.685 3.880 5.915 4.590 ;
        RECT 7.725 3.880 7.955 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 8.830 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.830 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.375 0.450 1.605 1.165 ;
        RECT 5.685 0.450 5.915 1.160 ;
        RECT 7.925 0.450 8.155 1.160 ;
        RECT 0.000 -0.450 8.400 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.255 2.060 0.585 3.685 ;
        RECT 2.925 3.505 4.890 3.685 ;
        RECT 2.925 3.455 6.355 3.505 ;
        RECT 2.925 2.875 3.155 3.455 ;
        RECT 4.665 3.275 6.355 3.455 ;
        RECT 2.320 2.415 3.715 2.645 ;
        RECT 2.320 2.060 2.550 2.415 ;
        RECT 3.945 2.185 4.175 3.215 ;
        RECT 0.255 1.830 2.550 2.060 ;
        RECT 3.155 1.955 4.175 2.185 ;
        RECT 0.255 0.845 0.485 1.830 ;
        RECT 3.155 1.490 3.385 1.955 ;
        RECT 4.665 1.655 4.895 3.275 ;
        RECT 6.125 2.450 6.355 3.275 ;
        RECT 2.495 1.085 3.385 1.490 ;
        RECT 3.615 1.315 4.895 1.655 ;
        RECT 5.125 1.825 6.410 2.055 ;
        RECT 5.125 1.085 5.355 1.825 ;
        RECT 2.495 0.680 5.355 1.085 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_2
MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.640 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.870 2.330 2.090 2.710 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.547000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 1.750 6.115 2.150 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.995200 ;
    PORT
      LAYER Metal1 ;
        RECT 7.895 3.140 8.125 3.720 ;
        RECT 9.935 3.140 10.165 3.720 ;
        RECT 7.895 2.910 10.165 3.140 ;
        RECT 9.045 1.650 9.390 2.910 ;
        RECT 7.865 1.390 10.335 1.650 ;
        RECT 7.865 0.840 8.095 1.390 ;
        RECT 10.105 0.840 10.335 1.390 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 10.640 5.490 ;
        RECT 1.365 3.845 1.595 4.590 ;
        RECT 4.655 4.035 4.885 4.590 ;
        RECT 6.695 3.565 6.925 4.590 ;
        RECT 8.915 3.880 9.145 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 11.070 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 11.070 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.165 ;
        RECT 4.270 0.450 4.610 0.680 ;
        RECT 6.510 0.450 6.850 0.680 ;
        RECT 8.985 0.450 9.215 1.160 ;
        RECT 0.000 -0.450 10.640 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.060 0.575 3.685 ;
        RECT 2.915 3.510 5.905 3.740 ;
        RECT 2.915 2.930 3.145 3.510 ;
        RECT 2.320 2.470 3.650 2.700 ;
        RECT 2.320 2.060 2.550 2.470 ;
        RECT 3.935 2.060 4.165 3.215 ;
        RECT 5.675 2.695 5.905 3.510 ;
        RECT 0.245 1.830 2.550 2.060 ;
        RECT 3.090 1.830 4.165 2.060 ;
        RECT 5.290 2.465 7.665 2.695 ;
        RECT 0.245 0.845 0.475 1.830 ;
        RECT 3.090 1.490 3.320 1.830 ;
        RECT 5.290 1.600 5.520 2.465 ;
        RECT 2.485 1.140 3.320 1.490 ;
        RECT 3.550 1.370 5.520 1.600 ;
        RECT 6.345 1.825 7.665 2.055 ;
        RECT 6.345 1.140 6.575 1.825 ;
        RECT 2.485 0.910 6.575 1.140 ;
        RECT 2.485 0.680 2.715 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_3
MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.760 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.870 2.330 2.090 2.710 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.735 1.770 6.115 2.150 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.244800 ;
    PORT
      LAYER Metal1 ;
        RECT 7.785 3.200 8.015 3.780 ;
        RECT 9.825 3.200 10.055 3.780 ;
        RECT 7.785 2.970 10.055 3.200 ;
        RECT 8.960 1.620 9.420 2.970 ;
        RECT 7.685 1.390 10.155 1.620 ;
        RECT 7.685 0.680 7.915 1.390 ;
        RECT 9.925 0.680 10.155 1.390 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 11.760 5.490 ;
        RECT 1.365 3.845 1.595 4.590 ;
        RECT 4.725 4.350 4.955 4.590 ;
        RECT 6.765 3.880 6.995 4.590 ;
        RECT 8.805 3.880 9.035 4.590 ;
        RECT 10.845 3.880 11.075 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 12.190 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.190 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.165 ;
        RECT 4.270 0.450 4.610 0.635 ;
        RECT 6.510 0.450 6.850 0.635 ;
        RECT 8.805 0.450 9.035 1.160 ;
        RECT 11.045 0.450 11.275 1.160 ;
        RECT 0.000 -0.450 11.760 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.060 0.575 3.685 ;
        RECT 2.915 3.510 4.625 3.740 ;
        RECT 2.915 2.930 3.145 3.510 ;
        RECT 2.320 2.470 3.650 2.700 ;
        RECT 2.320 2.060 2.550 2.470 ;
        RECT 3.935 2.060 4.165 3.215 ;
        RECT 0.245 1.830 2.550 2.060 ;
        RECT 3.090 1.830 4.165 2.060 ;
        RECT 4.395 2.735 4.625 3.510 ;
        RECT 5.745 2.735 5.975 3.720 ;
        RECT 4.395 2.505 8.560 2.735 ;
        RECT 0.245 0.845 0.475 1.830 ;
        RECT 3.090 1.490 3.320 1.830 ;
        RECT 4.395 1.600 4.625 2.505 ;
        RECT 2.485 1.140 3.320 1.490 ;
        RECT 3.550 1.370 4.625 1.600 ;
        RECT 6.345 1.850 8.560 2.080 ;
        RECT 6.345 1.140 6.575 1.850 ;
        RECT 2.485 0.910 6.575 1.140 ;
        RECT 2.485 0.680 2.715 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_4
MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.150 1.530 2.710 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.768000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.175 1.770 8.810 2.150 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.489600 ;
    PORT
      LAYER Metal1 ;
        RECT 10.015 3.080 16.365 3.835 ;
        RECT 15.760 1.650 16.365 3.080 ;
        RECT 15.760 1.595 17.065 1.650 ;
        RECT 10.115 0.865 17.065 1.595 ;
        RECT 16.835 0.840 17.065 0.865 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 18.480 5.490 ;
        RECT 1.265 3.845 1.495 4.590 ;
        RECT 4.915 3.880 5.145 4.590 ;
        RECT 6.955 3.880 7.185 4.590 ;
        RECT 8.995 3.880 9.225 4.590 ;
        RECT 11.035 4.350 11.265 4.590 ;
        RECT 13.075 4.350 13.305 4.590 ;
        RECT 15.115 4.350 15.345 4.590 ;
        RECT 17.155 3.880 17.385 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 18.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.695 ;
        RECT 4.270 0.450 4.610 0.625 ;
        RECT 6.755 0.450 6.985 0.690 ;
        RECT 8.995 0.450 9.225 0.690 ;
        RECT 11.180 0.450 11.520 0.635 ;
        RECT 13.420 0.450 13.760 0.635 ;
        RECT 15.660 0.450 16.000 0.635 ;
        RECT 17.955 0.450 18.185 1.160 ;
        RECT 0.000 -0.450 18.480 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.925 3.915 4.635 4.145 ;
        RECT 0.245 1.545 0.475 3.685 ;
        RECT 2.925 3.335 3.155 3.915 ;
        RECT 1.805 2.470 3.650 2.700 ;
        RECT 1.805 1.545 2.035 2.470 ;
        RECT 3.945 2.240 4.175 3.685 ;
        RECT 0.245 1.315 2.035 1.545 ;
        RECT 3.145 2.010 4.175 2.240 ;
        RECT 4.405 3.250 4.635 3.915 ;
        RECT 7.975 3.250 8.205 3.830 ;
        RECT 4.405 3.140 8.205 3.250 ;
        RECT 4.405 2.910 9.665 3.140 ;
        RECT 3.145 1.490 3.375 2.010 ;
        RECT 4.405 1.780 4.635 2.910 ;
        RECT 9.435 2.750 9.665 2.910 ;
        RECT 9.435 2.410 14.895 2.750 ;
        RECT 2.485 1.085 3.375 1.490 ;
        RECT 3.605 1.550 4.635 1.780 ;
        RECT 9.435 1.825 14.325 2.150 ;
        RECT 3.605 1.315 3.835 1.550 ;
        RECT 9.435 1.490 9.665 1.825 ;
        RECT 5.635 1.260 9.665 1.490 ;
        RECT 5.635 1.085 5.865 1.260 ;
        RECT 2.485 0.855 5.865 1.085 ;
        RECT 2.485 0.680 2.715 0.855 ;
        RECT 7.875 0.680 8.105 1.260 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_8
MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.200 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.330 1.575 2.710 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 10.151999 ;
    PORT
      LAYER Metal1 ;
        RECT 6.040 1.770 11.050 2.150 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.734400 ;
    PORT
      LAYER Metal1 ;
        RECT 12.255 3.365 22.685 4.175 ;
        RECT 22.080 1.650 22.685 3.365 ;
        RECT 22.080 1.600 23.785 1.650 ;
        RECT 12.355 0.865 23.785 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 25.200 5.490 ;
        RECT 1.505 3.845 1.735 4.590 ;
        RECT 5.115 3.880 5.345 4.590 ;
        RECT 7.155 3.880 7.385 4.590 ;
        RECT 9.195 3.880 9.425 4.590 ;
        RECT 11.235 3.880 11.465 4.590 ;
        RECT 13.220 4.405 13.560 4.590 ;
        RECT 15.260 4.405 15.600 4.590 ;
        RECT 17.300 4.405 17.640 4.590 ;
        RECT 19.340 4.405 19.680 4.590 ;
        RECT 21.380 4.405 21.720 4.590 ;
        RECT 23.475 3.880 23.705 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 25.630 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 25.630 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.695 ;
        RECT 4.270 0.450 4.610 0.625 ;
        RECT 6.700 0.450 7.040 0.635 ;
        RECT 8.940 0.450 9.280 0.635 ;
        RECT 11.180 0.450 11.520 0.635 ;
        RECT 13.420 0.450 13.760 0.635 ;
        RECT 15.660 0.450 16.000 0.635 ;
        RECT 17.900 0.450 18.240 0.635 ;
        RECT 20.140 0.450 20.480 0.635 ;
        RECT 22.380 0.450 22.720 0.635 ;
        RECT 24.675 0.450 24.905 1.160 ;
        RECT 0.000 -0.450 25.200 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.485 3.170 0.715 3.750 ;
        RECT 2.925 3.675 3.155 4.255 ;
        RECT 2.925 3.445 4.635 3.675 ;
        RECT 4.405 3.360 4.635 3.445 ;
        RECT 10.215 3.360 10.445 3.940 ;
        RECT 0.485 2.940 3.595 3.170 ;
        RECT 1.805 1.600 2.035 2.940 ;
        RECT 3.365 2.415 3.595 2.940 ;
        RECT 3.945 2.185 4.175 3.215 ;
        RECT 0.190 1.370 2.035 1.600 ;
        RECT 3.145 1.955 4.175 2.185 ;
        RECT 4.405 3.140 10.445 3.360 ;
        RECT 4.405 2.910 11.695 3.140 ;
        RECT 3.145 1.490 3.375 1.955 ;
        RECT 4.405 1.655 4.635 2.910 ;
        RECT 11.465 2.790 11.695 2.910 ;
        RECT 11.465 2.450 21.210 2.790 ;
        RECT 2.485 1.085 3.375 1.490 ;
        RECT 3.605 1.315 4.635 1.655 ;
        RECT 11.675 1.830 21.035 2.150 ;
        RECT 11.675 1.490 11.905 1.830 ;
        RECT 5.635 1.260 11.905 1.490 ;
        RECT 5.635 1.085 8.105 1.260 ;
        RECT 2.485 0.865 8.105 1.085 ;
        RECT 2.485 0.855 5.865 0.865 ;
        RECT 2.485 0.680 2.715 0.855 ;
        RECT 7.875 0.680 8.105 0.865 ;
        RECT 10.115 0.680 10.345 1.260 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_12
MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 31.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.545 2.330 1.575 2.710 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 13.535999 ;
    PORT
      LAYER Metal1 ;
        RECT 5.300 2.150 12.125 2.710 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 12.979199 ;
    PORT
      LAYER Metal1 ;
        RECT 14.520 3.365 29.090 4.175 ;
        RECT 28.530 1.650 29.090 3.365 ;
        RECT 28.530 1.635 30.505 1.650 ;
        RECT 14.595 0.865 30.505 1.635 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 31.920 5.490 ;
        RECT 1.505 3.845 1.735 4.590 ;
        RECT 4.860 4.370 5.200 4.590 ;
        RECT 6.900 4.370 7.240 4.590 ;
        RECT 8.940 4.370 9.280 4.590 ;
        RECT 11.280 4.370 11.620 4.590 ;
        RECT 13.500 4.405 13.840 4.590 ;
        RECT 15.540 4.405 15.880 4.590 ;
        RECT 17.580 4.405 17.920 4.590 ;
        RECT 19.620 4.405 19.960 4.590 ;
        RECT 21.660 4.405 22.000 4.590 ;
        RECT 23.700 4.405 24.040 4.590 ;
        RECT 25.740 4.405 26.080 4.590 ;
        RECT 27.780 4.405 28.120 4.590 ;
        RECT 29.875 3.880 30.105 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 32.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 32.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.695 ;
        RECT 4.270 0.450 4.610 0.625 ;
        RECT 6.700 0.450 7.040 0.635 ;
        RECT 8.940 0.450 9.280 0.635 ;
        RECT 11.180 0.450 11.520 0.635 ;
        RECT 13.405 0.450 13.780 0.635 ;
        RECT 15.660 0.450 16.000 0.635 ;
        RECT 17.900 0.450 18.240 0.635 ;
        RECT 20.140 0.450 20.480 0.635 ;
        RECT 22.380 0.450 22.720 0.635 ;
        RECT 24.620 0.450 24.960 0.635 ;
        RECT 26.860 0.450 27.200 0.635 ;
        RECT 29.100 0.450 29.440 0.635 ;
        RECT 31.395 0.450 31.625 1.160 ;
        RECT 0.000 -0.450 31.920 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.485 3.170 0.715 3.750 ;
        RECT 2.925 3.445 12.700 4.140 ;
        RECT 4.405 3.330 12.700 3.445 ;
        RECT 0.485 2.940 3.595 3.170 ;
        RECT 1.805 1.600 2.035 2.940 ;
        RECT 3.365 2.415 3.595 2.940 ;
        RECT 3.945 2.185 4.175 3.215 ;
        RECT 0.190 1.370 2.035 1.600 ;
        RECT 3.145 1.955 4.175 2.185 ;
        RECT 3.145 1.490 3.375 1.955 ;
        RECT 4.405 1.655 4.635 3.330 ;
        RECT 12.355 2.755 12.700 3.330 ;
        RECT 12.355 2.470 27.620 2.755 ;
        RECT 2.485 1.085 3.375 1.490 ;
        RECT 3.605 1.315 4.635 1.655 ;
        RECT 13.855 1.865 27.775 2.160 ;
        RECT 13.855 1.650 14.145 1.865 ;
        RECT 5.635 1.085 14.145 1.650 ;
        RECT 2.485 0.865 14.145 1.085 ;
        RECT 2.485 0.855 5.865 0.865 ;
        RECT 2.485 0.680 2.715 0.855 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_16
MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.676500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.740 1.015 2.550 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.157200 ;
    PORT
      LAYER Metal1 ;
        RECT 2.565 1.590 2.895 3.775 ;
        RECT 2.390 1.210 2.895 1.590 ;
        RECT 2.665 0.710 2.895 1.210 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 3.360 5.490 ;
        RECT 1.365 3.240 1.595 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 3.790 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 3.790 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.050 ;
        RECT 0.000 -0.450 3.360 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.010 0.575 3.775 ;
        RECT 0.345 2.780 2.215 3.010 ;
        RECT 1.930 1.740 2.215 2.780 ;
        RECT 1.930 1.510 2.160 1.740 ;
        RECT 0.245 1.280 2.160 1.510 ;
        RECT 0.245 0.710 0.475 1.280 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.353000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 2.000 0.970 3.270 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.550600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.665 3.960 3.110 4.300 ;
        RECT 2.880 1.215 3.110 3.960 ;
        RECT 2.330 0.710 3.110 1.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 4.480 5.490 ;
        RECT 1.265 3.960 1.495 4.590 ;
        RECT 3.685 3.550 3.915 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.215 ;
        RECT 3.785 0.450 4.015 1.215 ;
        RECT 0.000 -0.450 4.480 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.730 0.475 4.360 ;
        RECT 0.245 3.500 1.600 3.730 ;
        RECT 1.370 2.500 1.600 3.500 ;
        RECT 1.370 2.270 2.650 2.500 ;
        RECT 1.370 1.770 1.600 2.270 ;
        RECT 0.245 1.540 1.600 1.770 ;
        RECT 0.245 0.875 0.475 1.540 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_2
MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.035000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.805 2.215 1.975 2.555 ;
        RECT 0.805 1.770 1.530 2.215 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.329000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.785 3.190 4.015 4.230 ;
        RECT 5.925 3.190 6.255 4.230 ;
        RECT 3.785 2.960 6.255 3.190 ;
        RECT 5.750 1.875 6.255 2.960 ;
        RECT 3.785 1.645 6.255 1.875 ;
        RECT 3.785 1.075 4.015 1.645 ;
        RECT 5.750 1.075 6.255 1.645 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.840 5.490 ;
        RECT 0.245 3.420 0.475 4.590 ;
        RECT 2.385 3.420 2.615 4.590 ;
        RECT 4.805 3.420 5.035 4.590 ;
        RECT 7.045 3.420 7.275 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 8.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.415 ;
        RECT 2.665 0.450 2.895 1.415 ;
        RECT 4.905 0.450 5.135 1.415 ;
        RECT 7.145 0.450 7.375 1.415 ;
        RECT 0.000 -0.450 7.840 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 3.190 1.595 4.230 ;
        RECT 1.365 2.960 2.435 3.190 ;
        RECT 2.205 2.555 2.435 2.960 ;
        RECT 2.205 2.215 4.745 2.555 ;
        RECT 2.205 1.360 2.435 2.215 ;
        RECT 1.310 1.130 2.435 1.360 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_3
MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.706000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.805 2.215 1.975 2.555 ;
        RECT 0.805 1.770 1.530 2.215 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.101200 ;
    PORT
      LAYER Metal1 ;
        RECT 3.785 3.320 4.015 4.360 ;
        RECT 5.925 3.320 6.155 4.360 ;
        RECT 3.785 3.090 6.155 3.320 ;
        RECT 5.750 1.875 6.155 3.090 ;
        RECT 5.750 1.675 6.255 1.875 ;
        RECT 3.785 1.445 6.255 1.675 ;
        RECT 3.785 0.875 4.015 1.445 ;
        RECT 5.750 0.875 6.255 1.445 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.840 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.805 3.550 5.035 4.590 ;
        RECT 7.045 3.550 7.275 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 8.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.215 ;
        RECT 2.665 0.450 2.895 1.215 ;
        RECT 4.905 0.450 5.135 1.215 ;
        RECT 7.145 0.450 7.375 1.215 ;
        RECT 0.000 -0.450 7.840 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 1.365 3.090 2.435 3.320 ;
        RECT 2.205 2.555 2.435 3.090 ;
        RECT 2.205 2.215 4.745 2.555 ;
        RECT 2.205 1.160 2.435 2.215 ;
        RECT 1.310 0.930 2.435 1.160 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_4
MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.412000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 2.215 4.205 2.650 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.202400 ;
    PORT
      LAYER Metal1 ;
        RECT 6.025 3.320 6.255 4.360 ;
        RECT 8.165 3.320 8.395 4.360 ;
        RECT 10.230 3.320 10.635 4.360 ;
        RECT 12.645 3.320 12.875 4.360 ;
        RECT 6.025 3.090 12.875 3.320 ;
        RECT 9.150 1.745 9.650 3.090 ;
        RECT 6.025 1.515 12.975 1.745 ;
        RECT 6.025 0.945 6.255 1.515 ;
        RECT 8.265 0.945 8.495 1.515 ;
        RECT 10.505 0.945 10.735 1.515 ;
        RECT 12.745 0.945 12.975 1.515 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.560 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.875 4.855 4.590 ;
        RECT 7.045 3.550 7.275 4.590 ;
        RECT 9.285 3.550 9.515 4.590 ;
        RECT 11.525 3.550 11.755 4.590 ;
        RECT 13.765 3.550 13.995 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.285 ;
        RECT 2.485 0.450 2.715 1.285 ;
        RECT 4.725 0.450 4.955 1.285 ;
        RECT 7.145 0.450 7.375 1.285 ;
        RECT 9.385 0.450 9.615 1.215 ;
        RECT 11.625 0.450 11.855 1.215 ;
        RECT 13.865 0.450 14.095 1.285 ;
        RECT 0.000 -0.450 14.560 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 1.365 3.090 4.665 3.320 ;
        RECT 4.435 2.650 4.665 3.090 ;
        RECT 4.435 2.270 8.920 2.650 ;
        RECT 9.880 2.270 13.510 2.650 ;
        RECT 4.435 1.745 4.665 2.270 ;
        RECT 1.365 1.515 4.665 1.745 ;
        RECT 1.365 0.945 1.595 1.515 ;
        RECT 3.605 0.945 3.835 1.515 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_8
MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 8.118000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.275 2.215 6.675 2.555 ;
        RECT 1.275 1.770 6.010 2.215 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.303599 ;
    PORT
      LAYER Metal1 ;
        RECT 8.485 3.320 8.715 4.360 ;
        RECT 10.625 3.320 10.855 4.360 ;
        RECT 12.865 3.320 13.095 4.360 ;
        RECT 14.710 3.320 15.335 4.360 ;
        RECT 17.345 3.320 17.575 4.360 ;
        RECT 19.585 3.320 19.815 4.360 ;
        RECT 8.485 3.090 19.815 3.320 ;
        RECT 13.465 1.540 14.350 3.090 ;
        RECT 8.485 1.310 19.915 1.540 ;
        RECT 8.485 1.180 8.715 1.310 ;
        RECT 10.725 0.740 10.955 1.310 ;
        RECT 12.965 0.740 13.195 1.310 ;
        RECT 15.205 0.740 15.435 1.310 ;
        RECT 17.445 0.740 17.675 1.310 ;
        RECT 19.685 1.180 19.915 1.310 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 21.280 5.490 ;
        RECT 0.465 3.550 0.695 4.590 ;
        RECT 2.605 3.550 2.835 4.590 ;
        RECT 4.845 3.550 5.075 4.590 ;
        RECT 7.365 3.875 7.595 4.590 ;
        RECT 9.505 3.550 9.735 4.590 ;
        RECT 11.745 3.550 11.975 4.590 ;
        RECT 13.985 3.550 14.215 4.590 ;
        RECT 16.225 3.550 16.455 4.590 ;
        RECT 18.465 3.550 18.695 4.590 ;
        RECT 20.705 3.550 20.935 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 21.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.315 ;
        RECT 2.705 0.450 2.935 1.080 ;
        RECT 4.945 0.450 5.175 1.080 ;
        RECT 7.185 0.450 7.415 1.080 ;
        RECT 9.605 0.450 9.835 1.080 ;
        RECT 11.845 0.450 12.075 1.080 ;
        RECT 14.085 0.450 14.315 1.080 ;
        RECT 16.325 0.450 16.555 1.080 ;
        RECT 18.565 0.450 18.795 1.080 ;
        RECT 20.805 0.450 21.035 1.080 ;
        RECT 0.000 -0.450 21.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.585 3.320 1.815 4.360 ;
        RECT 3.725 3.320 3.955 4.360 ;
        RECT 5.965 3.320 6.195 4.360 ;
        RECT 1.585 3.090 7.135 3.320 ;
        RECT 6.905 2.555 7.135 3.090 ;
        RECT 6.905 2.215 13.205 2.555 ;
        RECT 14.580 2.215 19.980 2.555 ;
        RECT 6.905 1.540 7.135 2.215 ;
        RECT 1.585 1.310 7.135 1.540 ;
        RECT 1.585 1.110 1.815 1.310 ;
        RECT 3.825 1.110 4.055 1.310 ;
        RECT 6.065 1.110 6.295 1.310 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_12
MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.000 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 10.823999 ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 2.125 7.965 2.840 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 12.404799 ;
    PORT
      LAYER Metal1 ;
        RECT 10.505 3.320 10.735 4.360 ;
        RECT 12.645 3.320 12.875 4.360 ;
        RECT 14.885 3.320 15.115 4.360 ;
        RECT 17.125 3.320 17.355 4.360 ;
        RECT 19.365 3.320 19.595 4.360 ;
        RECT 21.605 3.320 21.835 4.360 ;
        RECT 23.845 3.320 24.075 4.360 ;
        RECT 26.085 3.320 26.315 4.360 ;
        RECT 10.505 3.090 26.315 3.320 ;
        RECT 17.985 1.895 18.735 3.090 ;
        RECT 10.505 1.745 18.735 1.895 ;
        RECT 10.505 1.665 26.415 1.745 ;
        RECT 10.505 1.515 12.975 1.665 ;
        RECT 10.505 0.945 10.735 1.515 ;
        RECT 12.745 0.945 12.975 1.515 ;
        RECT 14.985 0.945 15.215 1.665 ;
        RECT 17.225 1.515 26.415 1.665 ;
        RECT 17.225 0.945 17.455 1.515 ;
        RECT 19.465 0.945 19.695 1.515 ;
        RECT 21.705 0.945 21.935 1.515 ;
        RECT 23.945 0.945 24.175 1.515 ;
        RECT 26.185 0.945 26.415 1.515 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 28.000 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.875 9.335 4.590 ;
        RECT 11.525 3.550 11.755 4.590 ;
        RECT 13.765 3.550 13.995 4.590 ;
        RECT 16.005 3.550 16.235 4.590 ;
        RECT 18.245 3.550 18.475 4.590 ;
        RECT 20.485 3.550 20.715 4.590 ;
        RECT 22.725 3.550 22.955 4.590 ;
        RECT 24.965 3.550 25.195 4.590 ;
        RECT 27.205 3.550 27.435 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 28.430 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 28.430 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.285 ;
        RECT 2.485 0.450 2.715 1.285 ;
        RECT 4.725 0.450 4.955 1.285 ;
        RECT 6.965 0.450 7.195 1.285 ;
        RECT 9.205 0.450 9.435 1.285 ;
        RECT 11.625 0.450 11.855 1.285 ;
        RECT 13.865 0.450 14.095 1.285 ;
        RECT 16.105 0.450 16.335 1.215 ;
        RECT 18.345 0.450 18.575 1.215 ;
        RECT 20.585 0.450 20.815 1.285 ;
        RECT 22.825 0.450 23.055 1.215 ;
        RECT 25.065 0.450 25.295 1.215 ;
        RECT 27.305 0.450 27.535 1.285 ;
        RECT 0.000 -0.450 28.000 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 5.745 3.320 5.975 4.360 ;
        RECT 8.085 3.320 8.550 4.360 ;
        RECT 1.365 3.090 8.550 3.320 ;
        RECT 8.320 2.555 8.550 3.090 ;
        RECT 8.320 2.215 17.105 2.555 ;
        RECT 18.965 2.215 26.245 2.555 ;
        RECT 8.320 1.745 8.550 2.215 ;
        RECT 1.365 1.515 8.550 1.745 ;
        RECT 1.365 0.945 1.595 1.515 ;
        RECT 3.605 0.945 3.835 1.515 ;
        RECT 5.845 0.945 6.075 1.515 ;
        RECT 8.085 0.945 8.550 1.515 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_16
MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 ;
  ORIGIN 0.000 0.000 ;
  SIZE 34.720 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 13.530000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 2.215 9.845 2.650 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 15.506000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.745 3.320 12.975 4.360 ;
        RECT 14.885 3.320 15.115 4.360 ;
        RECT 17.125 3.320 17.355 4.360 ;
        RECT 19.365 3.320 19.595 4.360 ;
        RECT 21.605 3.320 21.835 4.360 ;
        RECT 23.845 3.320 24.075 4.360 ;
        RECT 26.085 3.320 26.315 4.360 ;
        RECT 28.325 3.320 28.555 4.360 ;
        RECT 30.565 3.320 30.795 4.360 ;
        RECT 32.805 3.320 33.035 4.360 ;
        RECT 12.745 3.090 33.035 3.320 ;
        RECT 22.465 1.745 23.215 3.090 ;
        RECT 12.745 1.675 23.215 1.745 ;
        RECT 12.745 1.515 33.135 1.675 ;
        RECT 12.745 0.945 13.005 1.515 ;
        RECT 14.985 0.945 15.215 1.515 ;
        RECT 17.225 0.945 17.455 1.515 ;
        RECT 19.465 0.945 19.695 1.515 ;
        RECT 21.705 1.445 33.135 1.515 ;
        RECT 21.705 0.945 21.935 1.445 ;
        RECT 23.945 0.945 24.175 1.445 ;
        RECT 26.185 0.945 26.415 1.445 ;
        RECT 28.425 0.945 28.655 1.445 ;
        RECT 30.665 0.945 30.895 1.445 ;
        RECT 32.905 0.945 33.135 1.445 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 34.720 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
        RECT 11.345 3.875 11.575 4.590 ;
        RECT 13.765 3.550 13.995 4.590 ;
        RECT 16.005 3.550 16.235 4.590 ;
        RECT 18.245 3.550 18.475 4.590 ;
        RECT 20.485 3.550 20.715 4.590 ;
        RECT 22.725 3.550 22.955 4.590 ;
        RECT 24.965 3.550 25.195 4.590 ;
        RECT 27.205 3.550 27.435 4.590 ;
        RECT 29.445 3.550 29.675 4.590 ;
        RECT 31.685 3.550 31.915 4.590 ;
        RECT 33.925 3.550 34.155 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 35.150 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 35.150 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.285 ;
        RECT 2.485 0.450 2.715 1.285 ;
        RECT 4.725 0.450 4.955 1.285 ;
        RECT 6.965 0.450 7.195 1.285 ;
        RECT 9.205 0.450 9.435 1.285 ;
        RECT 11.445 0.450 11.675 1.285 ;
        RECT 13.865 0.450 14.095 1.285 ;
        RECT 16.105 0.450 16.335 1.285 ;
        RECT 18.345 0.450 18.575 1.285 ;
        RECT 20.585 0.450 20.815 1.215 ;
        RECT 22.825 0.450 23.055 1.215 ;
        RECT 25.065 0.450 25.295 1.215 ;
        RECT 27.305 0.450 27.535 1.215 ;
        RECT 29.545 0.450 29.775 1.215 ;
        RECT 31.785 0.450 32.015 1.215 ;
        RECT 34.025 0.450 34.255 1.285 ;
        RECT 0.000 -0.450 34.720 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 5.745 3.320 5.975 4.360 ;
        RECT 7.985 3.320 8.215 4.360 ;
        RECT 10.225 3.320 10.455 4.360 ;
        RECT 1.365 3.090 10.455 3.320 ;
        RECT 10.225 2.650 10.455 3.090 ;
        RECT 10.225 2.215 21.225 2.650 ;
        RECT 23.445 2.215 32.605 2.650 ;
        RECT 10.225 1.745 10.555 2.215 ;
        RECT 1.365 1.515 10.555 1.745 ;
        RECT 1.365 0.945 1.595 1.515 ;
        RECT 3.605 0.945 3.835 1.515 ;
        RECT 5.845 0.945 6.075 1.515 ;
        RECT 8.085 0.945 8.315 1.515 ;
        RECT 10.325 0.945 10.555 1.515 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_20
MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.353000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 1.830 0.970 2.530 ;
        RECT 0.710 1.210 0.970 1.830 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.126400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 0.945 1.595 4.360 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 2.240 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 2.670 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.285 ;
        RECT 0.000 -0.450 2.240 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_1
MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.706000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.360 2.270 1.640 2.710 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.514200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.830 1.595 4.360 ;
        RECT 1.365 3.550 2.100 3.830 ;
        RECT 1.830 2.890 2.100 3.550 ;
        RECT 1.870 2.040 2.100 2.890 ;
        RECT 1.365 1.810 2.100 2.040 ;
        RECT 1.365 0.945 1.595 1.810 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 3.360 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 3.790 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 3.790 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.285 ;
        RECT 2.485 0.450 2.715 1.285 ;
        RECT 0.000 -0.450 3.360 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_2
MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.059000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 2.215 2.325 2.710 ;
        RECT 1.830 1.770 2.090 2.215 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.640600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.835 4.360 ;
        RECT 1.365 3.090 3.835 3.320 ;
        RECT 3.510 1.440 3.835 3.090 ;
        RECT 1.365 1.210 3.835 1.440 ;
        RECT 1.365 0.680 1.595 1.210 ;
        RECT 3.605 0.680 3.835 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 4.480 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.020 ;
        RECT 2.485 0.450 2.715 0.980 ;
        RECT 0.000 -0.450 4.480 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_3
MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.412000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 2.270 2.380 2.650 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.028400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.500 3.320 3.835 4.360 ;
        RECT 1.365 3.090 3.835 3.320 ;
        RECT 2.950 1.745 3.835 3.090 ;
        RECT 1.365 1.515 3.835 1.745 ;
        RECT 1.365 0.945 1.595 1.515 ;
        RECT 3.600 0.945 3.835 1.515 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.600 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.285 ;
        RECT 2.485 0.450 2.715 1.285 ;
        RECT 4.725 0.450 4.955 1.285 ;
        RECT 0.000 -0.450 5.600 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_4
MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 10.823999 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 2.265 4.260 2.645 ;
        RECT 5.360 2.215 8.880 2.650 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.056800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 5.745 3.320 5.975 4.360 ;
        RECT 7.985 3.320 8.215 4.360 ;
        RECT 1.365 3.090 8.215 3.320 ;
        RECT 4.630 1.745 5.130 3.090 ;
        RECT 1.365 1.515 8.315 1.745 ;
        RECT 1.365 0.945 1.625 1.515 ;
        RECT 3.605 0.945 3.835 1.515 ;
        RECT 5.845 0.945 6.075 1.515 ;
        RECT 8.085 0.945 8.315 1.515 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 10.080 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 10.510 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.285 ;
        RECT 2.485 0.450 2.715 1.285 ;
        RECT 4.725 0.450 4.955 1.285 ;
        RECT 6.965 0.450 7.195 1.285 ;
        RECT 9.205 0.450 9.435 1.285 ;
        RECT 0.000 -0.450 10.080 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_8
MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 16.236000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 2.270 6.140 2.650 ;
        RECT 7.660 2.270 13.170 2.650 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.085199 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 5.745 3.320 5.975 4.360 ;
        RECT 7.985 3.320 8.215 4.360 ;
        RECT 10.225 3.320 10.455 4.360 ;
        RECT 12.465 3.320 12.695 4.360 ;
        RECT 1.365 3.090 12.695 3.320 ;
        RECT 6.370 1.745 7.120 3.090 ;
        RECT 1.365 1.515 12.795 1.745 ;
        RECT 1.365 0.945 1.595 1.515 ;
        RECT 3.605 0.945 3.835 1.515 ;
        RECT 5.845 0.945 6.075 1.515 ;
        RECT 8.085 0.945 8.315 1.515 ;
        RECT 10.325 0.945 10.555 1.515 ;
        RECT 12.565 0.945 12.795 1.515 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.560 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
        RECT 11.345 3.550 11.575 4.590 ;
        RECT 13.585 3.550 13.815 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.285 ;
        RECT 2.485 0.450 2.715 1.285 ;
        RECT 4.725 0.450 4.955 1.285 ;
        RECT 6.965 0.450 7.195 1.285 ;
        RECT 9.205 0.450 9.435 1.285 ;
        RECT 11.445 0.450 11.675 1.285 ;
        RECT 13.685 0.450 13.915 1.285 ;
        RECT 0.000 -0.450 14.560 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_12
MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 21.647999 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 2.270 8.020 2.650 ;
        RECT 9.295 2.270 16.685 2.650 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 12.113600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 5.745 3.320 5.975 4.360 ;
        RECT 7.985 3.320 8.215 4.360 ;
        RECT 10.225 3.320 10.455 4.360 ;
        RECT 12.465 3.320 12.695 4.360 ;
        RECT 14.705 3.320 14.935 4.360 ;
        RECT 16.945 3.320 17.175 4.360 ;
        RECT 1.365 3.090 17.175 3.320 ;
        RECT 8.265 1.745 9.065 3.090 ;
        RECT 1.365 1.515 17.275 1.745 ;
        RECT 1.365 0.945 1.625 1.515 ;
        RECT 3.605 0.945 3.835 1.515 ;
        RECT 5.845 0.945 6.075 1.515 ;
        RECT 8.085 0.945 8.315 1.515 ;
        RECT 10.325 0.945 10.555 1.515 ;
        RECT 12.565 0.945 12.795 1.515 ;
        RECT 14.805 0.945 15.035 1.515 ;
        RECT 17.045 0.945 17.275 1.515 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 19.040 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
        RECT 11.345 3.550 11.575 4.590 ;
        RECT 13.585 3.550 13.815 4.590 ;
        RECT 15.825 3.550 16.055 4.590 ;
        RECT 18.065 3.550 18.295 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 19.470 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 19.470 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.285 ;
        RECT 2.485 0.450 2.715 1.285 ;
        RECT 4.725 0.450 4.955 1.285 ;
        RECT 6.965 0.450 7.195 1.285 ;
        RECT 9.205 0.450 9.435 1.285 ;
        RECT 11.445 0.450 11.675 1.285 ;
        RECT 13.685 0.450 13.915 1.285 ;
        RECT 15.925 0.450 16.155 1.285 ;
        RECT 18.165 0.450 18.395 1.285 ;
        RECT 0.000 -0.450 19.040 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_16
MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_20 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 27.059999 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 2.270 9.900 2.650 ;
        RECT 11.110 2.270 20.380 2.650 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 15.141999 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 5.745 3.320 5.975 4.360 ;
        RECT 7.985 3.320 8.215 4.360 ;
        RECT 10.225 3.320 10.455 4.360 ;
        RECT 12.465 3.320 12.695 4.360 ;
        RECT 14.705 3.320 14.935 4.360 ;
        RECT 16.945 3.320 17.175 4.360 ;
        RECT 19.185 3.320 19.415 4.360 ;
        RECT 21.425 3.320 21.655 4.360 ;
        RECT 1.365 3.090 21.655 3.320 ;
        RECT 10.130 1.745 10.880 3.090 ;
        RECT 1.365 1.515 21.755 1.745 ;
        RECT 1.365 0.945 1.625 1.515 ;
        RECT 3.605 0.945 3.835 1.515 ;
        RECT 5.845 0.945 6.075 1.515 ;
        RECT 8.085 0.945 8.315 1.515 ;
        RECT 10.325 0.945 10.555 1.515 ;
        RECT 12.565 0.945 12.795 1.515 ;
        RECT 14.805 0.945 15.035 1.515 ;
        RECT 17.045 0.945 17.275 1.515 ;
        RECT 19.285 0.945 19.515 1.515 ;
        RECT 21.525 0.945 21.755 1.515 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 23.520 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
        RECT 11.345 3.550 11.575 4.590 ;
        RECT 13.585 3.550 13.815 4.590 ;
        RECT 15.825 3.550 16.055 4.590 ;
        RECT 18.065 3.550 18.295 4.590 ;
        RECT 20.305 3.550 20.535 4.590 ;
        RECT 22.545 3.550 22.775 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 23.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 23.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.285 ;
        RECT 2.485 0.450 2.715 1.285 ;
        RECT 4.725 0.450 4.955 1.285 ;
        RECT 6.965 0.450 7.195 1.285 ;
        RECT 9.205 0.450 9.435 1.285 ;
        RECT 11.445 0.450 11.675 1.285 ;
        RECT 13.685 0.450 13.915 1.285 ;
        RECT 15.925 0.450 16.155 1.285 ;
        RECT 18.165 0.450 18.395 1.285 ;
        RECT 20.405 0.450 20.635 1.285 ;
        RECT 22.645 0.450 22.875 1.285 ;
        RECT 0.000 -0.450 23.520 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_20
MACRO gf180mcu_fd_sc_mcu9t5v0__dffnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.800 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 2.330 4.330 2.710 ;
    END
  END D
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.235 1.570 2.710 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.710 1.315 15.055 3.215 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 16.800 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.305 3.610 3.535 4.590 ;
        RECT 7.405 3.140 7.635 4.590 ;
        RECT 12.545 3.905 12.775 4.590 ;
        RECT 15.845 3.875 16.075 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 17.230 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 17.230 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.205 0.450 3.435 1.130 ;
        RECT 7.625 0.450 7.855 0.625 ;
        RECT 12.765 0.450 12.995 0.625 ;
        RECT 15.945 0.450 16.175 1.165 ;
        RECT 0.000 -0.450 16.800 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.765 4.125 6.170 4.355 ;
        RECT 0.345 3.170 0.575 3.750 ;
        RECT 3.765 3.220 3.995 4.125 ;
        RECT 0.345 2.940 2.035 3.170 ;
        RECT 1.805 1.740 2.035 2.940 ;
        RECT 0.245 1.510 2.035 1.740 ;
        RECT 2.385 2.990 3.995 3.220 ;
        RECT 0.245 1.315 0.475 1.510 ;
        RECT 2.385 1.315 2.715 2.990 ;
        RECT 4.425 2.970 4.790 3.780 ;
        RECT 4.560 1.360 4.790 2.970 ;
        RECT 4.325 1.020 4.790 1.360 ;
        RECT 5.445 2.280 5.675 3.780 ;
        RECT 8.965 2.850 9.195 3.780 ;
        RECT 6.965 2.510 9.195 2.850 ;
        RECT 5.445 2.050 8.515 2.280 ;
        RECT 5.445 1.020 5.675 2.050 ;
        RECT 8.285 1.940 8.515 2.050 ;
        RECT 6.125 1.085 6.355 1.820 ;
        RECT 8.965 1.315 9.195 2.510 ;
        RECT 10.085 2.990 10.315 3.780 ;
        RECT 11.470 3.445 15.515 3.675 ;
        RECT 10.085 2.760 13.410 2.990 ;
        RECT 10.085 1.315 10.315 2.760 ;
        RECT 10.545 2.300 11.250 2.530 ;
        RECT 13.925 2.460 14.155 3.215 ;
        RECT 12.050 2.455 14.155 2.460 ;
        RECT 10.545 1.085 10.775 2.300 ;
        RECT 12.050 2.230 14.480 2.455 ;
        RECT 14.105 1.315 14.480 2.230 ;
        RECT 6.125 0.855 10.775 1.085 ;
        RECT 11.425 1.085 11.655 1.225 ;
        RECT 15.285 1.085 15.515 3.445 ;
        RECT 11.425 0.855 15.515 1.085 ;
        RECT 9.350 0.680 10.775 0.855 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnq_1
MACRO gf180mcu_fd_sc_mcu9t5v0__dffnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.360 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 1.690 4.325 2.235 ;
    END
  END D
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.330 1.865 2.710 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.820 1.600 16.090 3.270 ;
        RECT 15.710 1.370 16.090 1.600 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.360 5.490 ;
        RECT 1.655 3.425 1.885 4.590 ;
        RECT 3.495 3.615 3.725 4.590 ;
        RECT 7.925 3.145 8.155 4.590 ;
        RECT 12.805 4.345 13.035 4.590 ;
        RECT 14.800 4.345 15.030 4.590 ;
        RECT 16.840 3.875 17.070 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 17.790 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 17.790 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.555 0.450 1.785 1.225 ;
        RECT 3.395 0.450 3.625 1.190 ;
        RECT 7.925 0.450 8.155 1.190 ;
        RECT 12.805 0.450 13.035 1.165 ;
        RECT 14.590 0.450 14.930 0.640 ;
        RECT 16.885 0.450 17.115 1.165 ;
        RECT 0.000 -0.450 17.360 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.955 4.130 6.690 4.360 ;
        RECT 0.635 3.170 0.865 3.750 ;
        RECT 3.955 3.215 4.185 4.130 ;
        RECT 0.635 2.940 2.325 3.170 ;
        RECT 2.095 1.740 2.325 2.940 ;
        RECT 0.435 1.510 2.325 1.740 ;
        RECT 2.675 2.985 4.185 3.215 ;
        RECT 0.435 1.315 0.665 1.510 ;
        RECT 2.675 1.315 2.905 2.985 ;
        RECT 4.515 2.975 4.790 3.785 ;
        RECT 4.560 1.080 4.790 2.975 ;
        RECT 5.965 2.285 6.195 3.785 ;
        RECT 8.945 2.855 9.175 3.785 ;
        RECT 7.485 2.625 9.175 2.855 ;
        RECT 7.485 2.515 7.715 2.625 ;
        RECT 8.365 2.285 8.595 2.395 ;
        RECT 5.965 2.055 8.595 2.285 ;
        RECT 8.945 2.285 9.175 2.625 ;
        RECT 10.385 2.880 10.615 3.785 ;
        RECT 11.785 3.690 16.550 3.920 ;
        RECT 11.785 3.110 12.015 3.690 ;
        RECT 10.385 2.650 13.530 2.880 ;
        RECT 8.945 2.055 9.495 2.285 ;
        RECT 5.965 1.080 6.195 2.055 ;
        RECT 6.590 1.595 9.035 1.825 ;
        RECT 8.805 0.910 9.035 1.595 ;
        RECT 9.265 1.315 9.495 2.055 ;
        RECT 10.385 1.315 10.615 2.650 ;
        RECT 13.190 2.470 13.530 2.650 ;
        RECT 11.170 2.190 11.550 2.420 ;
        RECT 11.170 0.910 11.400 2.190 ;
        RECT 13.825 2.150 14.055 3.215 ;
        RECT 12.310 2.060 14.055 2.150 ;
        RECT 12.310 1.920 15.525 2.060 ;
        RECT 13.870 1.830 15.525 1.920 ;
        RECT 11.630 1.395 13.640 1.625 ;
        RECT 11.630 1.370 11.970 1.395 ;
        RECT 13.410 1.140 13.640 1.395 ;
        RECT 13.870 1.370 14.210 1.830 ;
        RECT 16.320 1.140 16.550 3.690 ;
        RECT 13.410 0.910 16.550 1.140 ;
        RECT 8.805 0.680 11.400 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnq_2
MACRO gf180mcu_fd_sc_mcu9t5v0__dffnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.430 2.330 4.330 2.710 ;
    END
  END D
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.330 1.705 2.710 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.710 2.890 18.290 3.230 ;
        RECT 17.785 1.640 18.290 2.890 ;
        RECT 15.710 1.370 18.290 1.640 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 19.600 5.490 ;
        RECT 1.495 3.425 1.725 4.590 ;
        RECT 3.435 3.515 3.665 4.590 ;
        RECT 7.535 3.045 7.765 4.590 ;
        RECT 12.805 4.345 13.035 4.590 ;
        RECT 14.745 4.345 14.975 4.590 ;
        RECT 16.785 4.345 17.015 4.590 ;
        RECT 18.825 4.345 19.055 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 20.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 20.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.495 0.450 1.725 1.225 ;
        RECT 3.335 0.450 3.565 1.145 ;
        RECT 7.755 0.450 7.985 0.625 ;
        RECT 12.750 0.450 13.090 0.640 ;
        RECT 14.590 0.450 14.930 0.640 ;
        RECT 16.830 0.450 17.170 0.640 ;
        RECT 19.125 0.450 19.355 1.165 ;
        RECT 0.000 -0.450 19.600 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.895 4.030 6.300 4.260 ;
        RECT 0.475 3.170 0.705 3.750 ;
        RECT 3.895 3.215 4.125 4.030 ;
        RECT 0.475 2.940 2.165 3.170 ;
        RECT 1.935 2.005 2.165 2.940 ;
        RECT 0.375 1.775 2.165 2.005 ;
        RECT 2.515 2.985 4.125 3.215 ;
        RECT 0.375 1.315 0.605 1.775 ;
        RECT 2.515 1.315 2.845 2.985 ;
        RECT 4.555 2.875 4.790 3.685 ;
        RECT 4.560 1.375 4.790 2.875 ;
        RECT 4.455 1.035 4.790 1.375 ;
        RECT 5.575 2.240 5.805 3.685 ;
        RECT 9.030 2.700 9.265 3.685 ;
        RECT 7.040 2.470 9.265 2.700 ;
        RECT 5.575 2.010 8.585 2.240 ;
        RECT 5.575 1.035 5.805 2.010 ;
        RECT 8.355 1.900 8.585 2.010 ;
        RECT 6.200 1.085 6.540 1.780 ;
        RECT 9.035 1.315 9.265 2.470 ;
        RECT 10.155 3.215 10.385 3.685 ;
        RECT 11.730 3.500 18.750 3.730 ;
        RECT 10.155 2.985 11.855 3.215 ;
        RECT 10.155 1.315 10.385 2.985 ;
        RECT 11.165 1.085 11.395 2.755 ;
        RECT 11.625 2.700 11.855 2.985 ;
        RECT 11.625 2.470 13.530 2.700 ;
        RECT 13.825 2.210 14.055 3.215 ;
        RECT 13.825 2.150 17.555 2.210 ;
        RECT 12.310 1.920 17.555 2.150 ;
        RECT 13.870 1.870 17.555 1.920 ;
        RECT 6.200 0.855 11.395 1.085 ;
        RECT 9.420 0.680 11.395 0.855 ;
        RECT 11.685 1.140 11.915 1.490 ;
        RECT 13.870 1.370 14.210 1.870 ;
        RECT 18.520 1.140 18.750 3.500 ;
        RECT 11.685 0.910 18.750 1.140 ;
        RECT 11.685 0.680 11.915 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnq_4
MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.945 2.310 3.770 2.710 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.030000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.590 1.210 13.910 2.025 ;
    END
  END RN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.665 2.235 1.575 2.710 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.830 3.450 16.390 3.830 ;
        RECT 16.160 0.845 16.390 3.450 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.920 5.490 ;
        RECT 1.305 3.425 1.535 4.590 ;
        RECT 3.045 3.515 3.275 4.590 ;
        RECT 7.125 3.515 7.355 4.590 ;
        RECT 8.865 3.355 9.095 4.590 ;
        RECT 13.185 4.260 13.525 4.590 ;
        RECT 15.280 3.735 15.510 4.590 ;
        RECT 17.180 3.875 17.410 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 18.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.205 0.450 3.435 1.225 ;
        RECT 8.245 0.450 8.475 1.225 ;
        RECT 13.020 0.450 13.250 1.225 ;
        RECT 17.280 0.450 17.510 1.165 ;
        RECT 0.000 -0.450 17.920 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.505 3.975 5.755 4.315 ;
        RECT 0.285 3.170 0.515 3.750 ;
        RECT 2.325 3.285 2.555 3.685 ;
        RECT 3.505 3.285 3.735 3.975 ;
        RECT 0.285 2.940 2.035 3.170 ;
        RECT 1.805 1.740 2.035 2.940 ;
        RECT 0.245 1.510 2.035 1.740 ;
        RECT 2.325 3.055 3.735 3.285 ;
        RECT 0.245 1.315 0.475 1.510 ;
        RECT 2.325 1.315 2.715 3.055 ;
        RECT 4.065 1.510 4.295 3.685 ;
        RECT 5.085 2.995 5.315 3.685 ;
        RECT 6.105 3.275 6.335 3.855 ;
        RECT 8.145 3.275 8.375 3.855 ;
        RECT 6.105 3.045 8.375 3.275 ;
        RECT 5.085 2.815 5.670 2.995 ;
        RECT 5.085 2.765 9.590 2.815 ;
        RECT 5.445 2.585 9.590 2.765 ;
        RECT 4.065 1.280 4.610 1.510 ;
        RECT 5.445 1.225 5.675 2.585 ;
        RECT 9.885 2.360 10.115 3.995 ;
        RECT 9.640 2.180 10.115 2.360 ;
        RECT 6.670 2.130 10.115 2.180 ;
        RECT 10.780 3.765 14.950 3.995 ;
        RECT 10.780 3.185 11.135 3.765 ;
        RECT 6.125 1.685 6.355 2.025 ;
        RECT 6.670 1.950 9.865 2.130 ;
        RECT 6.125 1.455 9.405 1.685 ;
        RECT 9.175 0.995 9.405 1.455 ;
        RECT 9.635 1.225 9.865 1.950 ;
        RECT 10.320 0.995 10.550 2.025 ;
        RECT 10.780 1.225 11.010 3.185 ;
        RECT 11.345 0.995 11.575 3.065 ;
        RECT 11.900 1.225 12.155 3.525 ;
        RECT 12.580 3.295 14.490 3.525 ;
        RECT 12.580 2.725 12.810 3.295 ;
        RECT 14.260 2.495 14.490 3.295 ;
        RECT 14.720 2.725 14.950 3.765 ;
        RECT 14.260 2.265 15.930 2.495 ;
        RECT 15.440 1.975 15.930 2.265 ;
        RECT 15.440 1.315 15.670 1.975 ;
        RECT 9.175 0.765 11.575 0.995 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1
MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.945 1.770 3.895 2.150 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.255000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.380 1.675 14.410 2.150 ;
    END
  END RN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 1.575 2.245 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 17.510 3.450 17.915 3.830 ;
        RECT 17.685 0.845 17.915 3.450 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 19.600 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.225 3.045 3.455 4.590 ;
        RECT 7.305 3.515 7.535 4.590 ;
        RECT 9.045 3.440 9.275 4.590 ;
        RECT 13.525 4.345 13.755 4.590 ;
        RECT 15.845 3.875 16.075 4.590 ;
        RECT 16.665 3.875 16.895 4.590 ;
        RECT 18.705 3.875 18.935 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 20.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 20.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.080 ;
        RECT 3.205 0.450 3.435 1.310 ;
        RECT 8.425 0.450 8.655 1.310 ;
        RECT 13.425 0.450 13.655 1.310 ;
        RECT 16.565 0.450 16.795 1.165 ;
        RECT 18.805 0.450 19.035 1.165 ;
        RECT 0.000 -0.450 19.600 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.685 4.030 5.990 4.260 ;
        RECT 0.345 3.105 0.575 3.685 ;
        RECT 0.345 2.875 2.035 3.105 ;
        RECT 1.805 1.540 2.035 2.875 ;
        RECT 0.245 1.310 2.035 1.540 ;
        RECT 2.385 2.815 2.615 3.685 ;
        RECT 3.685 2.815 3.915 4.030 ;
        RECT 2.385 2.585 3.915 2.815 ;
        RECT 0.245 1.190 0.475 1.310 ;
        RECT 2.385 1.190 2.715 2.585 ;
        RECT 4.245 1.310 4.555 3.685 ;
        RECT 5.265 2.690 5.495 3.685 ;
        RECT 6.285 3.150 6.515 3.730 ;
        RECT 8.325 3.150 8.555 3.730 ;
        RECT 6.285 2.920 8.555 3.150 ;
        RECT 5.265 2.460 9.770 2.690 ;
        RECT 5.265 1.310 5.675 2.460 ;
        RECT 10.065 2.230 10.295 4.080 ;
        RECT 6.070 1.825 6.580 2.055 ;
        RECT 6.810 2.000 10.295 2.230 ;
        RECT 11.185 3.850 15.495 4.080 ;
        RECT 11.185 3.270 11.420 3.850 ;
        RECT 6.350 1.770 6.580 1.825 ;
        RECT 6.350 1.540 9.835 1.770 ;
        RECT 9.605 1.080 9.835 1.540 ;
        RECT 10.065 1.310 10.295 2.000 ;
        RECT 10.525 1.080 10.755 2.110 ;
        RECT 11.185 1.310 11.415 3.270 ;
        RECT 11.645 1.080 11.875 3.150 ;
        RECT 12.285 1.310 12.535 3.610 ;
        RECT 14.545 2.610 14.775 3.215 ;
        RECT 12.810 2.380 15.035 2.610 ;
        RECT 15.265 2.415 15.495 3.850 ;
        RECT 14.805 2.185 15.035 2.380 ;
        RECT 14.805 1.955 17.390 2.185 ;
        RECT 15.845 1.830 17.390 1.955 ;
        RECT 9.605 0.850 11.875 1.080 ;
        RECT 15.845 0.845 16.075 1.830 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2
MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.945 2.330 3.895 2.710 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.255000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.105 1.590 14.335 2.050 ;
        RECT 14.105 1.210 14.410 1.590 ;
    END
  END RN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.235 1.575 2.710 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 17.685 3.295 17.915 3.685 ;
        RECT 19.725 3.295 20.175 3.685 ;
        RECT 17.685 2.875 20.175 3.295 ;
        RECT 19.715 1.655 20.175 2.875 ;
        RECT 17.685 1.395 20.175 1.655 ;
        RECT 17.685 0.845 17.915 1.395 ;
        RECT 19.750 0.815 20.175 1.395 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 21.840 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.225 3.615 3.455 4.590 ;
        RECT 7.305 3.615 7.535 4.590 ;
        RECT 9.045 3.380 9.275 4.590 ;
        RECT 13.525 4.345 13.755 4.590 ;
        RECT 15.845 3.875 16.075 4.590 ;
        RECT 16.665 3.875 16.895 4.590 ;
        RECT 18.705 3.875 18.935 4.590 ;
        RECT 20.745 3.875 20.975 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 22.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 22.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.205 0.450 3.435 1.250 ;
        RECT 8.725 0.450 8.955 1.250 ;
        RECT 13.425 0.450 13.655 1.250 ;
        RECT 16.565 0.450 16.795 1.165 ;
        RECT 18.805 0.450 19.035 1.165 ;
        RECT 21.045 0.450 21.275 1.165 ;
        RECT 0.000 -0.450 21.840 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.685 4.130 5.990 4.360 ;
        RECT 0.345 3.170 0.575 3.750 ;
        RECT 2.385 3.385 2.615 3.685 ;
        RECT 3.685 3.385 3.915 4.130 ;
        RECT 0.345 2.940 2.035 3.170 ;
        RECT 1.805 2.005 2.035 2.940 ;
        RECT 0.245 1.775 2.035 2.005 ;
        RECT 2.385 3.155 3.915 3.385 ;
        RECT 0.245 1.315 0.475 1.775 ;
        RECT 2.385 1.315 2.715 3.155 ;
        RECT 4.245 1.250 4.555 3.785 ;
        RECT 5.265 2.915 5.495 3.785 ;
        RECT 6.285 3.375 6.515 3.955 ;
        RECT 8.325 3.375 8.555 3.955 ;
        RECT 6.285 3.145 8.555 3.375 ;
        RECT 5.265 2.685 9.770 2.915 ;
        RECT 5.265 1.250 5.675 2.685 ;
        RECT 10.065 2.455 10.295 4.020 ;
        RECT 6.810 2.225 10.295 2.455 ;
        RECT 6.070 1.765 9.835 1.995 ;
        RECT 9.605 1.020 9.835 1.765 ;
        RECT 10.065 1.250 10.295 2.225 ;
        RECT 11.185 3.790 15.300 4.020 ;
        RECT 11.185 3.210 11.420 3.790 ;
        RECT 10.525 1.020 10.755 2.050 ;
        RECT 11.185 1.250 11.415 3.210 ;
        RECT 11.645 1.020 11.875 3.090 ;
        RECT 12.285 1.250 12.535 3.550 ;
        RECT 14.555 2.550 14.840 3.215 ;
        RECT 12.810 2.320 14.840 2.550 ;
        RECT 15.070 2.700 15.300 3.790 ;
        RECT 15.070 2.470 15.550 2.700 ;
        RECT 14.610 2.240 14.840 2.320 ;
        RECT 15.845 2.240 19.485 2.275 ;
        RECT 14.610 2.015 19.485 2.240 ;
        RECT 14.610 2.010 16.075 2.015 ;
        RECT 9.605 0.790 11.875 1.020 ;
        RECT 15.845 0.845 16.075 2.010 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4
MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.945 2.330 3.975 2.710 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.965 2.200 17.770 2.760 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.545 2.330 15.575 2.805 ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.235 1.575 2.710 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.705 1.655 20.010 3.685 ;
        RECT 19.685 0.845 20.010 1.655 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 21.280 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.305 3.515 3.535 4.590 ;
        RECT 7.605 4.375 7.835 4.590 ;
        RECT 10.805 4.375 11.035 4.590 ;
        RECT 14.850 3.950 15.190 4.590 ;
        RECT 16.890 3.950 17.230 4.590 ;
        RECT 18.985 3.425 19.215 4.590 ;
        RECT 20.725 3.875 20.955 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 21.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.205 0.450 3.435 1.425 ;
        RECT 8.945 0.450 9.175 1.425 ;
        RECT 16.945 0.450 17.175 1.225 ;
        RECT 20.805 0.450 21.035 1.165 ;
        RECT 0.000 -0.450 21.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.765 4.145 6.070 4.260 ;
        RECT 12.485 4.145 12.715 4.315 ;
        RECT 3.765 3.915 12.715 4.145 ;
        RECT 0.345 3.170 0.575 3.750 ;
        RECT 2.385 3.285 2.615 3.685 ;
        RECT 3.765 3.285 3.995 3.915 ;
        RECT 0.345 2.940 2.035 3.170 ;
        RECT 1.805 1.740 2.035 2.940 ;
        RECT 0.245 1.510 2.035 1.740 ;
        RECT 2.385 3.055 3.995 3.285 ;
        RECT 0.245 1.315 0.655 1.510 ;
        RECT 2.385 1.315 2.715 3.055 ;
        RECT 4.325 1.315 4.555 3.685 ;
        RECT 5.345 2.915 5.575 3.685 ;
        RECT 6.365 3.345 9.075 3.685 ;
        RECT 9.565 3.445 12.275 3.685 ;
        RECT 9.565 3.345 11.655 3.445 ;
        RECT 5.345 2.685 10.235 2.915 ;
        RECT 5.825 1.315 6.055 2.685 ;
        RECT 10.005 2.575 10.235 2.685 ;
        RECT 7.105 2.345 7.335 2.455 ;
        RECT 11.390 2.345 11.655 3.345 ;
        RECT 12.045 2.875 12.275 3.445 ;
        RECT 13.065 3.455 18.690 3.685 ;
        RECT 7.105 2.115 11.655 2.345 ;
        RECT 6.285 1.885 6.515 2.115 ;
        RECT 6.285 1.655 11.195 1.885 ;
        RECT 10.965 0.910 11.195 1.655 ;
        RECT 11.425 1.315 11.655 2.115 ;
        RECT 13.065 1.655 13.295 3.455 ;
        RECT 14.085 2.115 14.315 3.215 ;
        RECT 12.545 1.315 13.295 1.655 ;
        RECT 13.665 2.100 14.315 2.115 ;
        RECT 15.925 2.100 16.155 3.215 ;
        RECT 17.965 2.885 18.230 3.225 ;
        RECT 13.665 1.870 16.155 2.100 ;
        RECT 16.505 1.970 16.735 2.115 ;
        RECT 18.000 2.025 18.230 2.885 ;
        RECT 18.460 2.415 18.690 3.455 ;
        RECT 18.910 2.025 19.475 2.315 ;
        RECT 18.000 1.975 19.475 2.025 ;
        RECT 18.000 1.970 19.135 1.975 ;
        RECT 13.665 1.315 13.895 1.870 ;
        RECT 14.325 0.910 14.555 1.640 ;
        RECT 14.985 1.315 15.215 1.870 ;
        RECT 16.505 1.740 19.135 1.970 ;
        RECT 18.905 1.315 19.135 1.740 ;
        RECT 10.965 0.680 14.555 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1
MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.400 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.390 1.770 4.330 2.150 ;
        RECT 3.990 1.210 4.330 1.770 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.755 2.320 17.770 2.710 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.270 1.210 15.610 2.060 ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 1.580 2.150 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 20.670 0.845 21.130 3.830 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 22.400 5.490 ;
        RECT 1.470 3.425 1.700 4.590 ;
        RECT 3.210 3.595 3.440 4.590 ;
        RECT 7.690 4.480 7.920 4.590 ;
        RECT 10.830 4.480 11.060 4.590 ;
        RECT 14.775 3.960 15.115 4.590 ;
        RECT 16.815 3.960 17.155 4.590 ;
        RECT 18.910 3.905 19.140 4.590 ;
        RECT 19.650 3.875 19.880 4.590 ;
        RECT 21.690 3.875 21.920 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 22.830 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 22.830 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.415 0.450 1.755 1.045 ;
        RECT 3.440 0.450 3.670 1.425 ;
        RECT 8.875 0.450 9.215 1.370 ;
        RECT 16.870 0.450 17.100 1.225 ;
        RECT 19.550 0.450 19.780 1.165 ;
        RECT 21.790 0.450 22.020 1.165 ;
        RECT 0.000 -0.450 22.400 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.670 4.250 5.975 4.340 ;
        RECT 12.455 4.250 12.795 4.350 ;
        RECT 3.670 4.020 12.795 4.250 ;
        RECT 0.450 3.105 0.680 3.685 ;
        RECT 3.670 3.215 3.900 4.020 ;
        RECT 0.450 2.875 2.140 3.105 ;
        RECT 1.910 1.540 2.140 2.875 ;
        RECT 0.350 1.310 2.140 1.540 ;
        RECT 2.490 2.985 3.900 3.215 ;
        RECT 4.230 3.185 4.460 3.765 ;
        RECT 0.350 1.190 0.580 1.310 ;
        RECT 2.490 1.190 2.820 2.985 ;
        RECT 4.230 2.955 4.790 3.185 ;
        RECT 4.560 1.315 4.790 2.955 ;
        RECT 5.250 2.750 5.480 3.765 ;
        RECT 6.520 3.450 9.160 3.790 ;
        RECT 6.520 2.980 6.750 3.450 ;
        RECT 9.650 3.305 9.880 3.790 ;
        RECT 9.650 3.075 10.780 3.305 ;
        RECT 9.650 2.980 9.880 3.075 ;
        RECT 10.090 2.750 10.320 2.845 ;
        RECT 5.250 2.520 10.320 2.750 ;
        RECT 5.680 1.315 5.910 2.520 ;
        RECT 10.090 2.505 10.320 2.520 ;
        RECT 10.550 2.455 10.780 3.075 ;
        RECT 12.070 2.455 12.300 3.775 ;
        RECT 7.100 2.275 10.005 2.290 ;
        RECT 10.550 2.275 12.300 2.455 ;
        RECT 7.100 2.225 12.300 2.275 ;
        RECT 13.090 3.730 14.635 3.775 ;
        RECT 13.090 3.545 18.690 3.730 ;
        RECT 6.360 1.720 6.590 2.115 ;
        RECT 7.100 2.060 11.440 2.225 ;
        RECT 7.100 1.950 7.330 2.060 ;
        RECT 9.920 2.045 11.440 2.060 ;
        RECT 7.530 1.720 9.835 1.830 ;
        RECT 6.360 1.600 9.835 1.720 ;
        RECT 6.360 1.490 7.730 1.600 ;
        RECT 9.605 0.910 9.835 1.600 ;
        RECT 11.210 1.315 11.440 2.045 ;
        RECT 13.090 1.900 13.320 3.545 ;
        RECT 14.495 3.500 18.690 3.545 ;
        RECT 12.330 1.670 13.320 1.900 ;
        RECT 12.330 1.315 12.560 1.670 ;
        RECT 14.110 1.480 14.340 3.305 ;
        RECT 13.450 1.370 14.340 1.480 ;
        RECT 13.450 1.140 15.040 1.370 ;
        RECT 14.810 0.980 15.040 1.140 ;
        RECT 15.850 0.980 16.080 3.225 ;
        RECT 17.890 2.910 18.230 3.250 ;
        RECT 18.000 2.115 18.230 2.910 ;
        RECT 18.460 2.425 18.690 3.500 ;
        RECT 18.000 2.090 20.320 2.115 ;
        RECT 16.375 1.860 20.320 2.090 ;
        RECT 18.830 1.775 20.320 1.860 ;
        RECT 18.830 1.315 19.060 1.775 ;
        RECT 9.605 0.680 14.380 0.910 ;
        RECT 14.810 0.750 16.080 0.980 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2
MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.640 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.055 2.330 3.890 2.710 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.950 2.710 17.210 3.270 ;
        RECT 16.950 2.480 17.515 2.710 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.270 1.770 15.530 2.765 ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.295 1.570 2.710 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 20.590 3.105 20.820 3.685 ;
        RECT 22.630 3.105 23.060 3.685 ;
        RECT 20.590 2.875 23.060 3.105 ;
        RECT 22.665 1.655 23.060 2.875 ;
        RECT 20.590 1.395 23.060 1.655 ;
        RECT 20.590 0.845 20.820 1.395 ;
        RECT 22.550 0.815 23.060 1.395 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 24.640 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.205 3.515 3.435 4.590 ;
        RECT 7.465 4.490 7.695 4.590 ;
        RECT 10.665 4.490 10.895 4.590 ;
        RECT 14.695 3.960 15.035 4.590 ;
        RECT 16.735 3.960 17.075 4.590 ;
        RECT 18.830 3.435 19.060 4.590 ;
        RECT 19.570 3.875 19.800 4.590 ;
        RECT 21.610 3.875 21.840 4.590 ;
        RECT 23.650 3.875 23.880 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 25.070 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 25.070 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.205 0.450 3.435 1.425 ;
        RECT 8.405 0.450 8.635 1.425 ;
        RECT 16.790 0.450 17.020 1.225 ;
        RECT 19.470 0.450 19.700 1.165 ;
        RECT 21.710 0.450 21.940 1.165 ;
        RECT 23.950 0.450 24.180 1.165 ;
        RECT 0.000 -0.450 24.640 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.665 4.030 12.630 4.260 ;
        RECT 0.345 3.170 0.575 3.750 ;
        RECT 2.385 3.285 2.615 3.685 ;
        RECT 3.665 3.285 3.895 4.030 ;
        RECT 0.345 2.940 2.035 3.170 ;
        RECT 1.805 2.005 2.035 2.940 ;
        RECT 0.245 1.775 2.035 2.005 ;
        RECT 2.385 3.055 3.895 3.285 ;
        RECT 0.245 1.315 0.475 1.775 ;
        RECT 2.385 1.315 2.715 3.055 ;
        RECT 4.225 1.315 4.555 3.685 ;
        RECT 5.245 2.915 5.475 3.685 ;
        RECT 6.285 3.350 8.935 3.800 ;
        RECT 9.425 3.570 12.135 3.800 ;
        RECT 9.425 3.460 11.515 3.570 ;
        RECT 5.245 2.685 10.095 2.915 ;
        RECT 5.245 1.315 5.675 2.685 ;
        RECT 9.865 2.575 10.095 2.685 ;
        RECT 6.865 2.345 7.095 2.455 ;
        RECT 11.285 2.345 11.515 3.460 ;
        RECT 11.905 2.875 12.135 3.570 ;
        RECT 12.925 3.500 18.500 3.730 ;
        RECT 6.865 2.115 11.515 2.345 ;
        RECT 6.125 1.885 6.355 2.115 ;
        RECT 6.125 1.655 11.055 1.885 ;
        RECT 10.825 0.910 11.055 1.655 ;
        RECT 11.285 1.315 11.515 2.115 ;
        RECT 12.925 1.655 13.155 3.500 ;
        RECT 13.945 1.655 14.175 3.215 ;
        RECT 12.405 1.315 13.155 1.655 ;
        RECT 13.525 1.540 14.175 1.655 ;
        RECT 15.770 1.540 16.000 3.225 ;
        RECT 17.810 2.115 18.040 3.225 ;
        RECT 18.270 2.425 18.500 3.500 ;
        RECT 20.010 2.115 22.435 2.290 ;
        RECT 17.810 2.060 22.435 2.115 ;
        RECT 16.295 2.005 22.435 2.060 ;
        RECT 16.295 1.830 20.240 2.005 ;
        RECT 13.525 1.310 16.000 1.540 ;
        RECT 18.750 1.775 20.240 1.830 ;
        RECT 18.750 1.315 18.980 1.775 ;
        RECT 10.825 0.680 14.455 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4
MACRO gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.160 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 2.330 4.550 2.710 ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.150 2.265 14.975 2.710 ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 1.770 1.530 2.150 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 18.145 1.590 18.375 3.685 ;
        RECT 18.070 0.845 18.375 1.590 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 20.160 5.490 ;
        RECT 1.265 3.425 1.495 4.590 ;
        RECT 3.005 3.905 3.235 4.590 ;
        RECT 7.245 3.905 7.475 4.590 ;
        RECT 9.725 3.905 9.955 4.590 ;
        RECT 13.805 3.915 14.035 4.590 ;
        RECT 16.345 3.175 16.575 4.590 ;
        RECT 19.165 3.875 19.395 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 20.590 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 20.590 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.080 ;
        RECT 3.225 0.450 3.455 1.425 ;
        RECT 7.425 0.450 7.655 1.425 ;
        RECT 16.305 0.450 16.535 1.420 ;
        RECT 19.265 0.450 19.495 1.165 ;
        RECT 0.000 -0.450 20.160 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.105 0.475 3.685 ;
        RECT 2.285 3.675 2.515 3.685 ;
        RECT 5.650 3.675 5.990 4.260 ;
        RECT 11.305 3.675 11.535 4.315 ;
        RECT 14.130 3.685 16.115 3.705 ;
        RECT 2.285 3.445 11.535 3.675 ;
        RECT 11.885 3.475 16.115 3.685 ;
        RECT 11.885 3.455 14.225 3.475 ;
        RECT 0.245 2.875 2.035 3.105 ;
        RECT 1.805 1.540 2.035 2.875 ;
        RECT 0.245 1.310 2.035 1.540 ;
        RECT 0.245 1.170 0.475 1.310 ;
        RECT 2.285 1.170 2.715 3.445 ;
        RECT 3.050 2.985 4.530 3.215 ;
        RECT 3.050 2.100 3.280 2.985 ;
        RECT 3.050 1.870 3.915 2.100 ;
        RECT 3.685 1.655 3.915 1.870 ;
        RECT 5.265 2.060 5.495 3.215 ;
        RECT 8.485 2.700 8.715 3.215 ;
        RECT 10.865 2.700 11.095 3.215 ;
        RECT 6.530 2.470 11.095 2.700 ;
        RECT 5.265 1.830 8.190 2.060 ;
        RECT 3.685 1.315 4.575 1.655 ;
        RECT 5.265 1.315 5.695 1.830 ;
        RECT 9.425 1.315 9.655 2.470 ;
        RECT 11.885 2.005 12.115 3.455 ;
        RECT 15.105 3.215 15.335 3.245 ;
        RECT 13.085 2.985 15.335 3.215 ;
        RECT 13.085 2.875 13.920 2.985 ;
        RECT 15.105 2.905 15.335 2.985 ;
        RECT 10.725 1.775 12.115 2.005 ;
        RECT 10.725 1.315 10.955 1.775 ;
        RECT 13.690 1.545 13.920 2.875 ;
        RECT 15.885 2.730 16.115 3.475 ;
        RECT 15.885 2.500 17.070 2.730 ;
        RECT 17.365 2.315 17.595 3.715 ;
        RECT 17.365 2.270 17.915 2.315 ;
        RECT 15.685 1.975 17.915 2.270 ;
        RECT 15.685 1.930 17.655 1.975 ;
        RECT 11.845 1.205 13.920 1.545 ;
        RECT 17.425 1.315 17.655 1.930 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1
MACRO gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.830 1.960 4.890 2.190 ;
        RECT 4.630 1.770 4.890 1.960 ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.655 2.165 14.860 2.710 ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.235 1.575 2.710 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.120 0.845 19.450 3.685 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 21.280 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.305 3.580 3.535 4.590 ;
        RECT 7.305 3.110 7.535 4.590 ;
        RECT 9.365 3.110 9.595 4.590 ;
        RECT 13.745 3.970 13.975 4.590 ;
        RECT 16.345 3.210 16.575 4.590 ;
        RECT 18.100 3.875 18.330 4.590 ;
        RECT 20.140 3.875 20.370 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 21.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.150 0.450 3.490 1.270 ;
        RECT 7.405 0.450 7.635 1.325 ;
        RECT 16.245 0.450 16.475 1.420 ;
        RECT 18.100 0.450 18.330 1.165 ;
        RECT 20.340 0.450 20.570 1.165 ;
        RECT 0.000 -0.450 21.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.765 4.095 7.075 4.325 ;
        RECT 0.345 3.170 0.575 3.710 ;
        RECT 3.765 3.215 3.995 4.095 ;
        RECT 0.345 2.940 2.035 3.170 ;
        RECT 0.345 2.900 0.575 2.940 ;
        RECT 1.805 2.005 2.035 2.940 ;
        RECT 0.245 1.775 2.035 2.005 ;
        RECT 2.385 2.985 3.995 3.215 ;
        RECT 0.245 1.315 0.475 1.775 ;
        RECT 2.385 1.315 2.715 2.985 ;
        RECT 4.325 2.650 4.555 3.750 ;
        RECT 3.370 2.420 4.555 2.650 ;
        RECT 3.370 1.730 3.600 2.420 ;
        RECT 5.445 1.960 5.675 3.750 ;
        RECT 6.845 2.880 7.075 4.095 ;
        RECT 7.765 3.980 9.135 4.210 ;
        RECT 7.765 2.880 7.995 3.980 ;
        RECT 6.845 2.650 7.995 2.880 ;
        RECT 8.325 2.420 8.555 3.750 ;
        RECT 8.905 2.880 9.135 3.980 ;
        RECT 9.825 3.975 11.435 4.315 ;
        RECT 9.825 2.880 10.055 3.975 ;
        RECT 8.905 2.650 10.055 2.880 ;
        RECT 10.765 2.420 10.995 3.685 ;
        RECT 6.810 2.190 10.995 2.420 ;
        RECT 11.785 3.510 16.115 3.740 ;
        RECT 5.445 1.730 8.130 1.960 ;
        RECT 3.370 1.550 3.940 1.730 ;
        RECT 3.370 1.500 4.555 1.550 ;
        RECT 3.715 1.320 4.555 1.500 ;
        RECT 4.325 1.210 4.555 1.320 ;
        RECT 5.445 1.215 5.675 1.730 ;
        RECT 9.365 1.215 9.595 2.190 ;
        RECT 11.785 1.960 12.015 3.510 ;
        RECT 10.665 1.730 12.015 1.960 ;
        RECT 13.025 2.940 15.275 3.280 ;
        RECT 10.665 1.215 10.895 1.730 ;
        RECT 13.025 1.500 13.255 2.940 ;
        RECT 15.885 2.765 16.115 3.510 ;
        RECT 15.885 2.535 17.070 2.765 ;
        RECT 17.365 2.115 17.595 3.750 ;
        RECT 15.625 1.775 18.770 2.115 ;
        RECT 11.785 1.160 13.875 1.500 ;
        RECT 17.365 1.315 17.595 1.775 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2
MACRO gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 2.330 4.525 2.710 ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.710 2.150 15.530 2.710 ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.240 1.575 2.710 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.665 3.105 19.895 3.685 ;
        RECT 21.705 3.105 22.135 3.685 ;
        RECT 19.665 2.875 22.135 3.105 ;
        RECT 21.655 1.655 22.135 2.875 ;
        RECT 19.665 1.395 22.135 1.655 ;
        RECT 19.665 0.845 19.895 1.395 ;
        RECT 21.430 0.815 22.135 1.395 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 23.520 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.105 3.860 3.335 4.590 ;
        RECT 7.345 3.905 7.575 4.590 ;
        RECT 9.825 3.905 10.055 4.590 ;
        RECT 14.205 3.915 14.435 4.590 ;
        RECT 16.745 3.155 16.975 4.590 ;
        RECT 18.645 3.875 18.875 4.590 ;
        RECT 20.685 3.875 20.915 4.590 ;
        RECT 22.725 3.875 22.955 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 23.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 23.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.225 0.450 3.455 1.425 ;
        RECT 7.525 0.450 7.755 1.425 ;
        RECT 16.525 0.450 16.755 1.425 ;
        RECT 18.545 0.450 18.775 1.165 ;
        RECT 20.785 0.450 21.015 1.165 ;
        RECT 23.025 0.450 23.255 1.165 ;
        RECT 0.000 -0.450 23.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.170 0.575 3.750 ;
        RECT 5.805 3.720 6.035 4.360 ;
        RECT 2.385 3.630 2.615 3.685 ;
        RECT 3.520 3.675 6.035 3.720 ;
        RECT 11.565 3.675 11.795 4.315 ;
        RECT 3.520 3.630 11.795 3.675 ;
        RECT 2.385 3.490 11.795 3.630 ;
        RECT 2.385 3.400 3.705 3.490 ;
        RECT 5.895 3.445 11.795 3.490 ;
        RECT 12.145 3.455 16.515 3.685 ;
        RECT 0.345 2.940 2.035 3.170 ;
        RECT 1.805 1.685 2.035 2.940 ;
        RECT 0.245 1.455 2.035 1.685 ;
        RECT 0.245 1.315 0.475 1.455 ;
        RECT 2.385 1.315 2.715 3.400 ;
        RECT 4.290 3.170 4.630 3.205 ;
        RECT 3.050 2.940 4.630 3.170 ;
        RECT 3.050 2.100 3.280 2.940 ;
        RECT 3.050 1.870 4.575 2.100 ;
        RECT 4.345 1.315 4.575 1.870 ;
        RECT 5.365 2.060 5.595 3.260 ;
        RECT 8.585 2.745 8.815 3.215 ;
        RECT 11.125 2.745 11.355 3.215 ;
        RECT 6.630 2.515 11.355 2.745 ;
        RECT 5.365 1.830 8.290 2.060 ;
        RECT 5.365 1.315 5.795 1.830 ;
        RECT 9.825 1.315 10.055 2.515 ;
        RECT 12.145 2.005 12.375 3.455 ;
        RECT 13.485 2.995 15.790 3.225 ;
        RECT 13.485 2.875 14.335 2.995 ;
        RECT 11.125 1.775 12.375 2.005 ;
        RECT 11.125 1.315 11.355 1.775 ;
        RECT 14.105 1.545 14.335 2.875 ;
        RECT 16.285 2.710 16.515 3.455 ;
        RECT 16.285 2.480 17.470 2.710 ;
        RECT 17.765 2.320 17.995 3.695 ;
        RECT 17.765 2.115 21.425 2.320 ;
        RECT 16.085 1.960 21.425 2.115 ;
        RECT 16.085 1.775 18.055 1.960 ;
        RECT 12.245 1.205 14.335 1.545 ;
        RECT 17.825 1.315 18.055 1.775 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4
MACRO gf180mcu_fd_sc_mcu9t5v0__dffq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.680 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.630 1.210 4.890 2.115 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.235 1.575 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.710 2.330 15.115 3.685 ;
        RECT 14.885 0.845 15.115 2.330 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 15.680 5.490 ;
        RECT 1.365 3.895 1.595 4.590 ;
        RECT 3.185 3.905 3.415 4.590 ;
        RECT 7.205 3.045 7.435 4.590 ;
        RECT 12.025 3.145 12.255 4.590 ;
        RECT 13.765 3.875 13.995 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 16.110 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 16.110 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.205 0.450 3.435 1.435 ;
        RECT 7.295 0.450 7.525 0.625 ;
        RECT 11.925 0.450 12.155 1.265 ;
        RECT 13.765 0.450 13.995 1.165 ;
        RECT 0.000 -0.450 15.680 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.655 0.575 4.235 ;
        RECT 5.885 3.675 6.115 4.315 ;
        RECT 1.940 3.655 6.115 3.675 ;
        RECT 0.345 3.445 6.115 3.655 ;
        RECT 0.345 3.425 2.035 3.445 ;
        RECT 1.805 2.005 2.035 3.425 ;
        RECT 2.385 2.755 2.615 3.215 ;
        RECT 5.165 2.755 5.395 3.215 ;
        RECT 2.385 2.525 4.075 2.755 ;
        RECT 0.245 1.775 2.035 2.005 ;
        RECT 3.845 1.895 4.075 2.525 ;
        RECT 0.245 1.315 0.475 1.775 ;
        RECT 2.485 1.665 4.075 1.895 ;
        RECT 2.485 1.315 2.715 1.665 ;
        RECT 3.845 0.920 4.075 1.665 ;
        RECT 5.165 2.415 7.875 2.755 ;
        RECT 5.165 1.315 5.395 2.415 ;
        RECT 8.225 2.115 8.455 3.685 ;
        RECT 6.685 1.775 8.455 2.115 ;
        RECT 8.225 1.655 8.455 1.775 ;
        RECT 9.745 3.455 11.795 3.685 ;
        RECT 8.225 1.315 8.855 1.655 ;
        RECT 9.745 1.315 9.975 3.455 ;
        RECT 10.505 1.085 10.735 2.755 ;
        RECT 11.565 2.700 11.795 3.455 ;
        RECT 11.565 2.470 12.750 2.700 ;
        RECT 13.045 2.115 13.275 3.685 ;
        RECT 11.265 2.060 13.275 2.115 ;
        RECT 11.265 1.830 14.490 2.060 ;
        RECT 11.265 1.775 13.275 1.830 ;
        RECT 13.045 1.315 13.275 1.775 ;
        RECT 5.665 0.920 10.735 1.085 ;
        RECT 3.845 0.855 10.735 0.920 ;
        RECT 3.845 0.690 5.890 0.855 ;
        RECT 9.010 0.690 10.735 0.855 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffq_1
MACRO gf180mcu_fd_sc_mcu9t5v0__dffq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.800 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.630 1.210 5.080 2.050 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 1.770 1.490 2.150 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.995 1.590 15.325 3.685 ;
        RECT 14.710 1.210 15.325 1.590 ;
        RECT 15.095 0.845 15.325 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 16.800 5.490 ;
        RECT 1.210 3.950 1.550 4.590 ;
        RECT 3.395 3.885 3.625 4.590 ;
        RECT 7.235 3.090 7.465 4.590 ;
        RECT 12.235 3.875 12.465 4.590 ;
        RECT 13.975 3.875 14.205 4.590 ;
        RECT 16.015 3.875 16.245 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 17.230 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 17.230 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.665 1.595 1.080 ;
        RECT 1.365 0.450 3.425 0.665 ;
        RECT 7.555 0.450 7.785 0.545 ;
        RECT 12.135 0.450 12.365 1.160 ;
        RECT 13.975 0.450 14.205 1.165 ;
        RECT 16.215 0.450 16.445 1.165 ;
        RECT 0.000 -0.450 16.800 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.675 0.475 4.235 ;
        RECT 3.855 4.020 6.145 4.360 ;
        RECT 0.245 3.655 3.300 3.675 ;
        RECT 3.855 3.655 4.085 4.020 ;
        RECT 0.245 3.445 4.085 3.655 ;
        RECT 0.245 3.425 2.035 3.445 ;
        RECT 3.205 3.425 4.085 3.445 ;
        RECT 1.805 1.540 2.035 3.425 ;
        RECT 0.245 1.310 2.035 1.540 ;
        RECT 2.385 2.800 2.615 3.215 ;
        RECT 5.375 2.800 5.605 3.730 ;
        RECT 2.385 2.570 4.285 2.800 ;
        RECT 0.245 1.170 0.475 1.310 ;
        RECT 2.385 1.170 2.715 2.570 ;
        RECT 4.055 0.980 4.285 2.570 ;
        RECT 5.375 2.460 8.085 2.800 ;
        RECT 5.375 1.305 5.605 2.460 ;
        RECT 8.835 2.105 9.065 3.730 ;
        RECT 6.655 1.765 9.065 2.105 ;
        RECT 8.835 1.310 9.065 1.765 ;
        RECT 9.955 3.500 12.055 3.730 ;
        RECT 9.955 1.310 10.185 3.500 ;
        RECT 10.715 1.005 10.945 2.800 ;
        RECT 11.825 2.700 12.055 3.500 ;
        RECT 11.825 2.470 12.960 2.700 ;
        RECT 13.255 2.110 13.485 3.685 ;
        RECT 11.475 2.060 13.485 2.110 ;
        RECT 11.475 1.830 14.700 2.060 ;
        RECT 11.475 1.770 13.485 1.830 ;
        RECT 5.995 0.980 10.945 1.005 ;
        RECT 4.055 0.775 10.945 0.980 ;
        RECT 13.255 0.840 13.485 1.770 ;
        RECT 4.055 0.680 6.100 0.775 ;
        RECT 9.220 0.685 10.945 0.775 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffq_2
MACRO gf180mcu_fd_sc_mcu9t5v0__dffq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.630 1.210 4.890 2.115 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.235 1.505 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.125 3.105 15.355 3.685 ;
        RECT 17.165 3.105 17.770 3.685 ;
        RECT 15.125 2.875 17.770 3.105 ;
        RECT 17.115 1.655 17.770 2.875 ;
        RECT 15.285 1.395 17.770 1.655 ;
        RECT 15.285 0.845 15.515 1.395 ;
        RECT 17.510 0.815 17.770 1.395 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 19.600 5.490 ;
        RECT 1.310 3.950 1.650 4.590 ;
        RECT 3.185 3.905 3.415 4.590 ;
        RECT 7.125 3.045 7.355 4.590 ;
        RECT 12.065 3.875 12.295 4.590 ;
        RECT 14.105 3.875 14.335 4.590 ;
        RECT 16.145 3.875 16.375 4.590 ;
        RECT 18.185 3.875 18.415 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 20.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 20.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.205 0.450 3.435 1.435 ;
        RECT 7.290 0.450 7.520 0.625 ;
        RECT 11.925 0.450 12.155 1.165 ;
        RECT 14.165 0.450 14.395 1.165 ;
        RECT 16.405 0.450 16.635 1.165 ;
        RECT 18.645 0.450 18.875 1.165 ;
        RECT 0.000 -0.450 19.600 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.675 0.575 4.235 ;
        RECT 5.805 3.675 6.035 4.315 ;
        RECT 0.345 3.445 6.035 3.675 ;
        RECT 0.345 3.425 2.035 3.445 ;
        RECT 1.805 2.005 2.035 3.425 ;
        RECT 2.385 2.755 2.615 3.215 ;
        RECT 5.165 2.755 5.395 3.215 ;
        RECT 2.385 2.525 4.075 2.755 ;
        RECT 0.245 1.775 2.035 2.005 ;
        RECT 3.845 1.895 4.075 2.525 ;
        RECT 0.245 1.315 0.475 1.775 ;
        RECT 2.485 1.665 4.075 1.895 ;
        RECT 2.485 1.315 2.715 1.665 ;
        RECT 3.845 0.920 4.075 1.665 ;
        RECT 5.165 2.415 8.175 2.755 ;
        RECT 5.165 1.315 5.395 2.415 ;
        RECT 8.620 2.115 8.855 3.685 ;
        RECT 6.685 1.775 8.855 2.115 ;
        RECT 8.625 1.315 8.855 1.775 ;
        RECT 9.745 3.455 11.935 3.685 ;
        RECT 9.745 1.315 9.975 3.455 ;
        RECT 10.625 1.085 10.855 2.755 ;
        RECT 11.705 2.700 11.935 3.455 ;
        RECT 11.705 2.470 12.790 2.700 ;
        RECT 13.085 2.315 13.315 3.685 ;
        RECT 13.085 2.115 16.885 2.315 ;
        RECT 11.265 1.975 16.885 2.115 ;
        RECT 11.265 1.775 13.310 1.975 ;
        RECT 5.665 0.920 10.855 1.085 ;
        RECT 3.845 0.855 10.855 0.920 ;
        RECT 3.845 0.690 5.890 0.855 ;
        RECT 9.010 0.690 10.855 0.855 ;
        RECT 13.045 0.845 13.310 1.775 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffq_4
MACRO gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.280 2.330 3.915 2.710 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.830000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.865 1.660 14.380 2.000 ;
        RECT 14.150 1.590 14.380 1.660 ;
        RECT 14.150 1.210 15.070 1.590 ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.660 2.150 0.970 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.345 2.190 16.650 3.685 ;
        RECT 16.325 0.845 16.650 2.190 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.920 5.490 ;
        RECT 1.285 3.425 1.515 4.590 ;
        RECT 3.245 3.615 3.475 4.590 ;
        RECT 7.325 3.615 7.555 4.590 ;
        RECT 9.065 3.330 9.295 4.590 ;
        RECT 13.365 4.190 13.595 4.590 ;
        RECT 15.625 3.310 15.855 4.590 ;
        RECT 17.365 3.875 17.595 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 18.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.385 0.450 1.615 1.225 ;
        RECT 3.225 0.450 3.455 1.200 ;
        RECT 8.705 0.450 8.935 1.200 ;
        RECT 13.185 0.450 13.415 1.200 ;
        RECT 17.445 0.450 17.675 1.165 ;
        RECT 0.000 -0.450 17.920 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.705 4.130 4.990 4.360 ;
        RECT 0.265 3.170 0.495 3.685 ;
        RECT 2.305 3.385 2.535 3.685 ;
        RECT 3.705 3.385 3.935 4.130 ;
        RECT 0.265 2.940 1.430 3.170 ;
        RECT 0.265 2.875 0.495 2.940 ;
        RECT 1.200 2.260 1.430 2.940 ;
        RECT 2.305 3.155 3.935 3.385 ;
        RECT 1.200 2.030 2.010 2.260 ;
        RECT 1.200 1.685 1.430 2.030 ;
        RECT 0.210 1.455 1.430 1.685 ;
        RECT 0.210 1.370 1.085 1.455 ;
        RECT 2.305 1.315 2.735 3.155 ;
        RECT 4.265 1.200 4.575 3.785 ;
        RECT 5.285 2.915 5.515 3.785 ;
        RECT 6.305 3.375 6.535 3.955 ;
        RECT 8.345 3.375 8.575 3.955 ;
        RECT 6.305 3.145 8.575 3.375 ;
        RECT 5.285 2.685 9.790 2.915 ;
        RECT 5.285 1.540 5.520 2.685 ;
        RECT 10.085 2.460 10.315 3.970 ;
        RECT 9.855 2.405 10.315 2.460 ;
        RECT 6.830 2.230 10.315 2.405 ;
        RECT 10.945 3.960 11.335 3.970 ;
        RECT 10.945 3.730 15.295 3.960 ;
        RECT 10.945 3.160 11.335 3.730 ;
        RECT 6.830 2.175 10.055 2.230 ;
        RECT 5.850 1.715 9.595 1.945 ;
        RECT 5.285 1.200 5.695 1.540 ;
        RECT 9.365 0.970 9.595 1.715 ;
        RECT 9.825 1.200 10.055 2.175 ;
        RECT 10.285 0.970 10.515 2.000 ;
        RECT 10.945 1.200 11.175 3.160 ;
        RECT 11.485 0.970 11.830 2.985 ;
        RECT 12.065 1.200 12.355 3.500 ;
        RECT 14.605 2.650 14.835 3.500 ;
        RECT 15.065 2.700 15.295 3.730 ;
        RECT 12.650 2.470 14.835 2.650 ;
        RECT 12.650 2.240 16.100 2.470 ;
        RECT 15.605 1.290 15.835 2.240 ;
        RECT 9.365 0.740 11.830 0.970 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
MACRO gf180mcu_fd_sc_mcu9t5v0__dffrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.960 2.330 3.895 2.710 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.255000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.590 2.330 14.015 2.710 ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.265 1.590 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.601600 ;
    PORT
      LAYER Metal1 ;
        RECT 17.445 0.845 17.770 3.685 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 19.040 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.225 3.615 3.455 4.590 ;
        RECT 7.305 3.615 7.535 4.590 ;
        RECT 9.045 3.320 9.275 4.590 ;
        RECT 13.345 4.345 13.575 4.590 ;
        RECT 15.385 3.875 15.615 4.590 ;
        RECT 16.425 3.875 16.655 4.590 ;
        RECT 18.465 3.875 18.695 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 19.470 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 19.470 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.200 ;
        RECT 3.205 0.450 3.435 1.195 ;
        RECT 8.425 0.450 8.655 1.195 ;
        RECT 13.135 0.450 13.365 1.195 ;
        RECT 16.325 0.450 16.555 1.235 ;
        RECT 18.565 0.450 18.795 1.235 ;
        RECT 0.000 -0.450 19.040 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.685 4.130 4.970 4.360 ;
        RECT 0.345 3.195 0.575 3.735 ;
        RECT 2.385 3.385 2.615 3.685 ;
        RECT 3.685 3.385 3.915 4.130 ;
        RECT 0.345 2.965 2.090 3.195 ;
        RECT 0.345 2.925 0.575 2.965 ;
        RECT 1.860 2.035 2.090 2.965 ;
        RECT 0.245 1.805 2.090 2.035 ;
        RECT 2.385 3.155 3.915 3.385 ;
        RECT 0.245 1.290 0.475 1.805 ;
        RECT 2.385 1.290 2.715 3.155 ;
        RECT 4.245 1.195 4.555 3.785 ;
        RECT 5.265 2.915 5.495 3.785 ;
        RECT 6.285 3.375 6.515 3.955 ;
        RECT 8.325 3.375 8.555 3.955 ;
        RECT 6.285 3.145 8.555 3.375 ;
        RECT 5.265 2.685 9.770 2.915 ;
        RECT 5.265 1.525 5.495 2.685 ;
        RECT 10.065 2.455 10.295 3.960 ;
        RECT 6.810 2.225 10.295 2.455 ;
        RECT 10.895 3.730 15.155 3.960 ;
        RECT 5.855 1.710 9.535 1.940 ;
        RECT 5.265 1.185 5.675 1.525 ;
        RECT 9.305 0.965 9.535 1.710 ;
        RECT 9.765 1.195 9.995 2.225 ;
        RECT 10.225 0.965 10.455 1.995 ;
        RECT 10.895 1.195 11.315 3.730 ;
        RECT 11.555 2.690 11.815 3.030 ;
        RECT 11.555 0.965 11.785 2.690 ;
        RECT 12.105 1.535 12.335 3.490 ;
        RECT 12.630 2.940 14.695 3.170 ;
        RECT 12.630 2.745 12.970 2.940 ;
        RECT 14.465 2.185 14.695 2.940 ;
        RECT 14.925 2.415 15.155 3.730 ;
        RECT 14.465 1.955 17.050 2.185 ;
        RECT 12.015 1.195 12.335 1.535 ;
        RECT 15.555 1.830 17.050 1.955 ;
        RECT 9.305 0.735 11.785 0.965 ;
        RECT 15.555 0.725 15.785 1.830 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrnq_2
MACRO gf180mcu_fd_sc_mcu9t5v0__dffrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.890 1.750 3.895 2.090 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.123000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.970 1.750 13.780 2.090 ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.330 1.570 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 17.370 3.215 17.605 3.685 ;
        RECT 19.410 3.215 19.840 3.685 ;
        RECT 17.370 2.875 19.840 3.215 ;
        RECT 19.595 1.625 19.840 2.875 ;
        RECT 17.370 1.395 19.840 1.625 ;
        RECT 17.370 0.815 17.600 1.395 ;
        RECT 19.610 0.815 19.840 1.395 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 21.280 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.105 3.090 3.335 4.590 ;
        RECT 7.185 3.560 7.415 4.590 ;
        RECT 8.925 3.390 9.155 4.590 ;
        RECT 13.330 4.345 13.560 4.590 ;
        RECT 15.370 3.875 15.605 4.590 ;
        RECT 16.345 3.875 16.580 4.590 ;
        RECT 18.390 4.585 20.660 4.590 ;
        RECT 18.390 3.875 18.620 4.585 ;
        RECT 20.430 3.875 20.660 4.585 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 21.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.225 0.450 3.455 1.370 ;
        RECT 8.305 0.450 8.535 1.370 ;
        RECT 13.110 0.640 13.340 1.370 ;
        RECT 13.110 0.450 16.535 0.640 ;
        RECT 18.490 0.450 18.720 1.165 ;
        RECT 20.730 0.450 20.960 1.165 ;
        RECT 0.000 -0.450 21.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.665 4.020 4.795 4.360 ;
        RECT 0.345 3.170 0.575 3.750 ;
        RECT 0.345 2.940 2.035 3.170 ;
        RECT 1.805 1.685 2.035 2.940 ;
        RECT 0.245 1.455 2.035 1.685 ;
        RECT 2.385 2.860 2.615 3.685 ;
        RECT 3.665 2.860 3.895 4.020 ;
        RECT 2.385 2.630 3.895 2.860 ;
        RECT 2.385 1.600 2.615 2.630 ;
        RECT 0.245 1.315 0.475 1.455 ;
        RECT 2.385 1.260 2.715 1.600 ;
        RECT 4.125 1.260 4.575 3.730 ;
        RECT 5.145 2.860 5.375 3.730 ;
        RECT 6.165 3.320 6.395 3.900 ;
        RECT 8.205 3.320 8.435 3.900 ;
        RECT 6.165 3.090 8.435 3.320 ;
        RECT 5.145 2.630 9.650 2.860 ;
        RECT 5.145 1.600 5.375 2.630 ;
        RECT 9.995 2.430 10.225 4.030 ;
        RECT 9.765 2.290 10.225 2.430 ;
        RECT 6.690 2.200 10.225 2.290 ;
        RECT 10.870 3.800 15.060 4.030 ;
        RECT 10.870 3.220 11.245 3.800 ;
        RECT 6.690 2.060 9.980 2.200 ;
        RECT 6.145 1.830 6.375 2.060 ;
        RECT 6.145 1.600 9.520 1.830 ;
        RECT 5.145 1.260 5.695 1.600 ;
        RECT 9.290 1.030 9.520 1.600 ;
        RECT 9.750 1.260 9.980 2.060 ;
        RECT 10.410 1.030 10.640 2.060 ;
        RECT 10.870 1.260 11.100 3.220 ;
        RECT 11.455 1.030 11.685 3.100 ;
        RECT 11.990 1.260 12.265 3.560 ;
        RECT 12.670 2.760 14.580 3.215 ;
        RECT 14.350 2.185 14.580 2.760 ;
        RECT 14.830 2.415 15.060 3.800 ;
        RECT 14.350 1.955 19.365 2.185 ;
        RECT 15.530 1.315 15.760 1.955 ;
        RECT 9.290 0.800 11.685 1.030 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrnq_4
MACRO gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.720 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.965 2.545 3.770 2.710 ;
        RECT 2.965 2.315 4.010 2.545 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.300 2.330 17.210 2.890 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.710 2.890 15.055 3.270 ;
        RECT 14.825 2.470 15.055 2.890 ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.480 1.580 3.270 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.125 0.845 19.450 3.685 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 20.720 5.490 ;
        RECT 1.265 3.960 1.495 4.590 ;
        RECT 3.005 3.560 3.235 4.590 ;
        RECT 7.245 4.490 7.475 4.590 ;
        RECT 10.445 4.490 10.675 4.590 ;
        RECT 14.330 4.005 14.670 4.590 ;
        RECT 16.370 4.005 16.710 4.590 ;
        RECT 18.465 3.480 18.695 4.590 ;
        RECT 20.205 3.875 20.435 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 21.150 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.150 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.385 0.450 1.615 1.225 ;
        RECT 3.285 0.450 3.515 1.425 ;
        RECT 8.585 0.450 8.815 1.425 ;
        RECT 16.360 0.450 16.590 1.225 ;
        RECT 20.245 0.450 20.475 1.165 ;
        RECT 0.000 -0.450 20.720 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.465 4.020 4.835 4.360 ;
        RECT 5.570 4.260 5.910 4.305 ;
        RECT 5.570 4.030 12.490 4.260 ;
        RECT 0.245 3.500 2.055 3.730 ;
        RECT 0.245 3.390 0.475 3.500 ;
        RECT 1.825 1.740 2.055 3.500 ;
        RECT 0.265 1.510 2.055 1.740 ;
        RECT 2.285 3.330 2.515 3.750 ;
        RECT 3.465 3.330 3.695 4.020 ;
        RECT 2.285 3.100 3.695 3.330 ;
        RECT 0.265 1.315 0.495 1.510 ;
        RECT 2.285 1.315 2.735 3.100 ;
        RECT 4.025 3.005 4.255 3.730 ;
        RECT 4.025 2.775 4.635 3.005 ;
        RECT 4.405 1.315 4.635 2.775 ;
        RECT 5.045 2.915 5.275 3.730 ;
        RECT 6.065 3.350 8.715 3.800 ;
        RECT 9.205 3.570 11.855 3.800 ;
        RECT 9.205 3.460 9.955 3.570 ;
        RECT 5.045 2.685 9.495 2.915 ;
        RECT 5.525 1.315 5.755 2.685 ;
        RECT 9.265 2.575 9.495 2.685 ;
        RECT 6.805 2.345 7.035 2.455 ;
        RECT 9.725 2.345 9.955 3.460 ;
        RECT 11.625 2.875 11.855 3.570 ;
        RECT 12.645 3.545 18.135 3.775 ;
        RECT 12.645 3.195 12.875 3.545 ;
        RECT 12.085 2.965 12.875 3.195 ;
        RECT 12.085 2.645 12.315 2.965 ;
        RECT 13.665 2.735 13.895 3.215 ;
        RECT 11.665 2.415 12.315 2.645 ;
        RECT 12.785 2.505 14.495 2.735 ;
        RECT 6.805 2.115 10.775 2.345 ;
        RECT 5.985 1.885 6.215 2.115 ;
        RECT 5.985 1.655 10.315 1.885 ;
        RECT 10.085 0.910 10.315 1.655 ;
        RECT 10.545 1.315 10.775 2.115 ;
        RECT 11.665 1.315 11.895 2.415 ;
        RECT 12.785 1.315 13.015 2.505 ;
        RECT 13.295 0.910 13.525 2.275 ;
        RECT 14.265 2.240 14.495 2.505 ;
        RECT 15.405 2.240 15.635 3.270 ;
        RECT 14.265 2.010 15.635 2.240 ;
        RECT 17.445 2.060 17.675 3.270 ;
        RECT 17.905 2.470 18.135 3.545 ;
        RECT 18.320 2.060 18.895 2.315 ;
        RECT 14.265 1.315 14.630 2.010 ;
        RECT 15.865 1.975 18.895 2.060 ;
        RECT 15.865 1.830 18.550 1.975 ;
        RECT 18.320 1.315 18.550 1.830 ;
        RECT 10.085 0.680 13.525 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1
MACRO gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.945 2.500 3.770 2.710 ;
        RECT 2.945 2.270 4.010 2.500 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.040 2.330 17.275 2.710 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.220 1.770 15.115 2.150 ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 2.200 1.575 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 20.245 0.845 20.570 3.685 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 21.840 5.490 ;
        RECT 1.265 3.425 1.495 4.590 ;
        RECT 3.005 3.515 3.235 4.590 ;
        RECT 7.305 4.490 7.535 4.590 ;
        RECT 10.505 4.490 10.735 4.590 ;
        RECT 14.390 3.950 14.730 4.590 ;
        RECT 16.430 3.950 16.770 4.590 ;
        RECT 18.525 3.425 18.755 4.590 ;
        RECT 19.245 3.875 19.475 4.590 ;
        RECT 21.285 3.875 21.515 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 22.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 22.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.285 0.450 3.515 1.425 ;
        RECT 8.645 0.450 8.875 1.425 ;
        RECT 16.405 0.450 16.635 1.225 ;
        RECT 19.125 0.450 19.355 1.165 ;
        RECT 21.365 0.450 21.595 1.165 ;
        RECT 0.000 -0.450 21.840 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.465 3.975 4.835 4.315 ;
        RECT 5.570 4.030 12.550 4.260 ;
        RECT 0.245 3.170 0.475 3.750 ;
        RECT 2.285 3.285 2.515 3.685 ;
        RECT 3.465 3.285 3.695 3.975 ;
        RECT 0.245 2.940 2.035 3.170 ;
        RECT 1.805 1.740 2.035 2.940 ;
        RECT 0.245 1.510 2.035 1.740 ;
        RECT 2.285 3.055 3.695 3.285 ;
        RECT 0.245 1.315 0.475 1.510 ;
        RECT 2.285 1.315 2.715 3.055 ;
        RECT 4.025 2.960 4.255 3.685 ;
        RECT 5.045 3.105 5.275 3.685 ;
        RECT 6.065 3.350 8.775 3.800 ;
        RECT 9.265 3.570 11.915 3.800 ;
        RECT 9.265 3.460 10.835 3.570 ;
        RECT 4.025 2.730 4.635 2.960 ;
        RECT 5.045 2.875 9.555 3.105 ;
        RECT 4.405 1.315 4.635 2.730 ;
        RECT 5.525 1.315 5.755 2.875 ;
        RECT 9.325 2.575 9.555 2.875 ;
        RECT 6.805 2.345 7.035 2.455 ;
        RECT 10.605 2.345 10.835 3.460 ;
        RECT 11.685 2.875 11.915 3.570 ;
        RECT 12.705 3.455 18.195 3.685 ;
        RECT 6.805 2.115 10.835 2.345 ;
        RECT 5.985 1.885 6.215 2.115 ;
        RECT 5.985 1.655 10.375 1.885 ;
        RECT 10.145 0.910 10.375 1.655 ;
        RECT 10.605 1.315 10.835 2.115 ;
        RECT 12.705 2.110 12.935 3.455 ;
        RECT 11.725 1.880 12.935 2.110 ;
        RECT 11.725 1.315 11.955 1.880 ;
        RECT 13.725 1.650 13.955 3.215 ;
        RECT 12.845 1.540 13.955 1.650 ;
        RECT 15.450 2.875 15.695 3.215 ;
        RECT 15.450 1.540 15.680 2.875 ;
        RECT 17.505 2.115 17.735 3.215 ;
        RECT 17.965 2.415 18.195 3.455 ;
        RECT 17.505 2.100 19.795 2.115 ;
        RECT 15.910 1.870 19.795 2.100 ;
        RECT 12.845 1.200 15.680 1.540 ;
        RECT 18.365 1.775 19.795 1.870 ;
        RECT 18.365 1.315 18.595 1.775 ;
        RECT 10.145 0.680 13.790 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2
MACRO gf180mcu_fd_sc_mcu9t5v0__dffrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.080 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.945 2.500 3.770 2.710 ;
        RECT 2.945 2.270 4.010 2.500 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.185 2.330 17.275 2.710 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.260 1.770 15.115 2.150 ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 2.200 1.575 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 20.205 3.105 20.495 3.685 ;
        RECT 22.305 3.105 22.885 3.685 ;
        RECT 20.205 2.875 22.885 3.105 ;
        RECT 22.300 1.655 22.885 2.875 ;
        RECT 20.205 1.395 22.885 1.655 ;
        RECT 20.205 0.845 20.435 1.395 ;
        RECT 22.445 0.845 22.885 1.395 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 24.080 5.490 ;
        RECT 1.265 3.425 1.495 4.590 ;
        RECT 3.005 3.515 3.235 4.590 ;
        RECT 7.305 4.490 7.535 4.590 ;
        RECT 10.505 4.490 10.735 4.590 ;
        RECT 14.390 3.950 14.730 4.590 ;
        RECT 16.430 3.950 16.770 4.590 ;
        RECT 18.525 3.425 18.755 4.590 ;
        RECT 19.245 3.875 19.475 4.590 ;
        RECT 21.285 3.875 21.515 4.590 ;
        RECT 23.325 3.875 23.555 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 24.510 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 24.510 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.285 0.450 3.515 1.425 ;
        RECT 8.645 0.450 8.875 1.425 ;
        RECT 16.405 0.450 16.635 1.225 ;
        RECT 19.085 0.450 19.315 1.165 ;
        RECT 21.325 0.450 21.555 1.165 ;
        RECT 23.565 0.450 23.795 1.165 ;
        RECT 0.000 -0.450 24.080 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.465 3.975 4.835 4.315 ;
        RECT 5.570 4.030 12.550 4.260 ;
        RECT 0.245 3.170 0.475 3.750 ;
        RECT 2.285 3.285 2.515 3.685 ;
        RECT 3.465 3.285 3.695 3.975 ;
        RECT 0.245 2.940 2.035 3.170 ;
        RECT 1.805 1.740 2.035 2.940 ;
        RECT 0.245 1.510 2.035 1.740 ;
        RECT 2.285 3.055 3.695 3.285 ;
        RECT 0.245 1.315 0.475 1.510 ;
        RECT 2.285 1.315 2.715 3.055 ;
        RECT 4.025 2.960 4.255 3.685 ;
        RECT 5.045 3.105 5.275 3.685 ;
        RECT 6.065 3.350 8.775 3.800 ;
        RECT 9.265 3.570 11.915 3.800 ;
        RECT 9.265 3.460 10.835 3.570 ;
        RECT 4.025 2.730 4.635 2.960 ;
        RECT 5.045 2.875 9.555 3.105 ;
        RECT 4.405 1.315 4.635 2.730 ;
        RECT 5.525 1.315 5.755 2.875 ;
        RECT 9.325 2.575 9.555 2.875 ;
        RECT 6.805 2.345 7.035 2.455 ;
        RECT 10.605 2.345 10.835 3.460 ;
        RECT 11.685 2.875 11.915 3.570 ;
        RECT 12.705 3.455 18.195 3.685 ;
        RECT 6.805 2.115 10.835 2.345 ;
        RECT 5.985 1.885 6.215 2.115 ;
        RECT 5.985 1.655 10.375 1.885 ;
        RECT 10.145 0.910 10.375 1.655 ;
        RECT 10.605 1.315 10.835 2.115 ;
        RECT 12.705 2.110 12.935 3.455 ;
        RECT 11.725 1.880 12.935 2.110 ;
        RECT 11.725 1.315 11.955 1.880 ;
        RECT 13.725 1.650 13.955 3.215 ;
        RECT 12.845 1.540 13.955 1.650 ;
        RECT 15.450 2.875 15.695 3.215 ;
        RECT 15.450 1.540 15.680 2.875 ;
        RECT 17.505 2.115 17.735 3.215 ;
        RECT 17.965 2.415 18.195 3.455 ;
        RECT 19.520 2.115 22.070 2.315 ;
        RECT 17.505 2.100 22.070 2.115 ;
        RECT 15.910 1.975 22.070 2.100 ;
        RECT 15.910 1.870 19.755 1.975 ;
        RECT 12.845 1.200 15.680 1.540 ;
        RECT 18.365 1.865 19.755 1.870 ;
        RECT 18.365 1.315 18.595 1.865 ;
        RECT 10.145 0.680 13.790 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrsnq_4
MACRO gf180mcu_fd_sc_mcu9t5v0__dffsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.160 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 1.770 4.030 2.150 ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.970 1.830 14.655 2.170 ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.330 1.530 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.190 0.845 19.450 3.685 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 20.160 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.305 3.145 3.535 4.590 ;
        RECT 7.525 3.960 7.755 4.590 ;
        RECT 10.005 4.005 10.235 4.590 ;
        RECT 13.985 3.145 14.215 4.590 ;
        RECT 16.025 3.615 16.255 4.590 ;
        RECT 18.185 3.875 18.415 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 20.590 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 20.590 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.205 0.450 3.435 1.245 ;
        RECT 7.405 0.450 7.635 1.245 ;
        RECT 16.245 0.450 16.475 1.265 ;
        RECT 18.085 0.450 18.315 1.165 ;
        RECT 0.000 -0.450 20.160 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.765 4.130 5.150 4.360 ;
        RECT 0.345 3.170 0.575 3.750 ;
        RECT 0.345 2.940 2.035 3.170 ;
        RECT 1.805 2.005 2.035 2.940 ;
        RECT 0.245 1.775 2.035 2.005 ;
        RECT 2.385 2.915 2.615 3.685 ;
        RECT 3.765 2.915 3.995 4.130 ;
        RECT 2.385 2.685 3.995 2.915 ;
        RECT 0.245 1.315 0.475 1.775 ;
        RECT 2.385 1.315 2.715 2.685 ;
        RECT 4.325 1.135 4.555 3.785 ;
        RECT 5.445 2.340 5.675 3.785 ;
        RECT 5.970 3.730 6.310 4.360 ;
        RECT 11.345 3.775 11.575 4.315 ;
        RECT 7.895 3.730 11.575 3.775 ;
        RECT 5.970 3.545 11.575 3.730 ;
        RECT 5.970 3.500 8.035 3.545 ;
        RECT 8.765 2.975 11.135 3.315 ;
        RECT 8.765 2.800 10.015 2.975 ;
        RECT 6.810 2.570 10.015 2.800 ;
        RECT 5.445 2.110 8.470 2.340 ;
        RECT 5.445 1.135 5.675 2.110 ;
        RECT 6.070 1.650 8.095 1.880 ;
        RECT 7.865 0.910 8.095 1.650 ;
        RECT 9.785 1.315 10.015 2.570 ;
        RECT 11.925 2.115 12.155 3.685 ;
        RECT 13.265 2.915 13.495 3.685 ;
        RECT 15.005 2.915 15.235 3.785 ;
        RECT 13.265 2.685 15.235 2.915 ;
        RECT 15.585 2.730 17.455 3.215 ;
        RECT 13.265 2.630 13.495 2.685 ;
        RECT 10.905 1.885 12.155 2.115 ;
        RECT 12.510 2.400 13.495 2.630 ;
        RECT 15.585 2.515 18.855 2.730 ;
        RECT 10.905 1.030 11.135 1.885 ;
        RECT 12.510 1.655 12.740 2.400 ;
        RECT 17.365 2.390 18.855 2.515 ;
        RECT 12.025 1.600 12.740 1.655 ;
        RECT 14.885 1.830 16.970 2.060 ;
        RECT 12.025 1.260 14.215 1.600 ;
        RECT 14.885 1.030 15.115 1.830 ;
        RECT 17.365 1.315 17.595 2.390 ;
        RECT 7.865 0.680 10.510 0.910 ;
        RECT 10.905 0.800 15.115 1.030 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffsnq_1
MACRO gf180mcu_fd_sc_mcu9t5v0__dffsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.720 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.075 1.770 3.975 2.150 ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.435 1.590 14.665 2.115 ;
        RECT 14.435 1.210 14.970 1.590 ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.240 1.390 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.125 0.845 19.450 3.685 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 20.720 5.490 ;
        RECT 1.365 3.895 1.595 4.590 ;
        RECT 3.305 3.615 3.535 4.590 ;
        RECT 7.475 3.615 7.705 4.590 ;
        RECT 9.875 3.830 10.105 4.590 ;
        RECT 13.855 3.515 14.085 4.590 ;
        RECT 15.895 3.045 16.125 4.590 ;
        RECT 18.105 3.875 18.335 4.590 ;
        RECT 20.145 3.875 20.375 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 21.150 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.150 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.205 0.450 3.435 1.320 ;
        RECT 7.475 0.450 7.705 1.320 ;
        RECT 16.115 0.450 16.345 1.165 ;
        RECT 18.005 0.450 18.235 1.165 ;
        RECT 20.245 0.450 20.475 1.165 ;
        RECT 0.000 -0.450 20.720 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.765 4.130 5.295 4.360 ;
        RECT 0.345 3.010 2.035 3.240 ;
        RECT 3.765 3.215 3.995 4.130 ;
        RECT 0.345 2.900 0.575 3.010 ;
        RECT 1.805 1.740 2.035 3.010 ;
        RECT 0.245 1.510 2.035 1.740 ;
        RECT 2.385 2.985 3.995 3.215 ;
        RECT 0.245 1.315 0.475 1.510 ;
        RECT 2.385 1.315 2.715 2.985 ;
        RECT 4.325 1.210 4.555 3.785 ;
        RECT 5.445 2.415 5.820 3.785 ;
        RECT 6.115 3.385 6.455 4.360 ;
        RECT 7.935 3.600 9.650 3.775 ;
        RECT 11.215 3.675 11.445 4.315 ;
        RECT 10.275 3.600 11.445 3.675 ;
        RECT 7.935 3.545 11.445 3.600 ;
        RECT 7.935 3.385 8.165 3.545 ;
        RECT 6.115 3.155 8.165 3.385 ;
        RECT 9.425 3.445 11.445 3.545 ;
        RECT 9.425 3.370 10.445 3.445 ;
        RECT 8.575 2.800 8.805 3.315 ;
        RECT 10.775 2.800 11.005 3.215 ;
        RECT 6.980 2.570 11.005 2.800 ;
        RECT 5.445 2.340 6.810 2.415 ;
        RECT 5.445 2.185 8.420 2.340 ;
        RECT 5.445 1.210 5.675 2.185 ;
        RECT 6.640 2.110 8.420 2.185 ;
        RECT 6.130 1.880 6.470 1.955 ;
        RECT 6.130 1.650 8.165 1.880 ;
        RECT 7.935 0.910 8.165 1.650 ;
        RECT 9.655 1.315 9.885 2.570 ;
        RECT 11.795 2.115 12.025 3.685 ;
        RECT 14.875 3.215 15.105 3.795 ;
        RECT 11.435 1.885 12.025 2.115 ;
        RECT 13.135 2.985 15.105 3.215 ;
        RECT 10.775 0.980 11.005 1.425 ;
        RECT 11.435 0.980 11.665 1.885 ;
        RECT 13.135 1.655 13.365 2.985 ;
        RECT 17.135 2.630 17.445 3.685 ;
        RECT 15.455 2.290 17.445 2.630 ;
        RECT 17.215 2.115 17.445 2.290 ;
        RECT 11.895 1.550 13.365 1.655 ;
        RECT 15.200 1.830 16.840 2.060 ;
        RECT 11.895 1.210 14.165 1.550 ;
        RECT 15.200 0.980 15.430 1.830 ;
        RECT 7.935 0.680 10.380 0.910 ;
        RECT 10.775 0.750 15.430 0.980 ;
        RECT 17.215 1.775 18.775 2.115 ;
        RECT 17.215 0.845 17.465 1.775 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffsnq_2
MACRO gf180mcu_fd_sc_mcu9t5v0__dffsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.945 2.330 4.030 2.710 ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.530 2.220 14.515 2.710 ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.240 1.570 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.110 3.105 19.340 3.685 ;
        RECT 21.150 3.105 21.880 3.685 ;
        RECT 19.110 2.875 21.880 3.105 ;
        RECT 21.590 1.655 21.880 2.875 ;
        RECT 19.405 1.395 21.880 1.655 ;
        RECT 19.405 0.845 19.640 1.395 ;
        RECT 21.590 0.845 21.880 1.395 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 23.520 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.305 3.615 3.535 4.590 ;
        RECT 7.510 3.615 7.740 4.590 ;
        RECT 9.715 3.885 10.055 4.590 ;
        RECT 13.790 3.515 14.020 4.590 ;
        RECT 15.830 3.045 16.060 4.590 ;
        RECT 18.090 3.875 18.320 4.590 ;
        RECT 20.130 3.875 20.360 4.590 ;
        RECT 22.170 3.875 22.400 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 23.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 23.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.225 ;
        RECT 3.205 0.450 3.435 1.425 ;
        RECT 7.455 0.450 7.795 1.370 ;
        RECT 15.995 0.450 16.335 0.640 ;
        RECT 18.290 0.450 18.520 1.165 ;
        RECT 20.530 0.450 20.760 1.165 ;
        RECT 22.770 0.450 23.000 1.165 ;
        RECT 0.000 -0.450 23.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.765 4.130 5.295 4.360 ;
        RECT 0.345 3.170 0.575 3.750 ;
        RECT 2.385 3.385 2.615 3.685 ;
        RECT 3.765 3.385 3.995 4.130 ;
        RECT 0.345 2.940 2.090 3.170 ;
        RECT 1.860 1.685 2.090 2.940 ;
        RECT 0.245 1.455 2.090 1.685 ;
        RECT 2.385 3.155 3.995 3.385 ;
        RECT 0.245 1.315 0.475 1.455 ;
        RECT 2.385 1.315 2.715 3.155 ;
        RECT 4.325 1.315 4.555 3.785 ;
        RECT 5.445 2.520 5.820 3.785 ;
        RECT 6.115 3.385 6.455 4.360 ;
        RECT 7.970 3.655 9.545 3.720 ;
        RECT 11.150 3.655 11.380 4.315 ;
        RECT 7.970 3.490 11.380 3.655 ;
        RECT 7.970 3.385 8.200 3.490 ;
        RECT 9.320 3.425 11.380 3.490 ;
        RECT 6.115 3.155 8.200 3.385 ;
        RECT 8.475 2.800 8.815 3.260 ;
        RECT 10.655 2.800 10.995 3.160 ;
        RECT 7.015 2.570 10.995 2.800 ;
        RECT 5.445 2.340 6.790 2.520 ;
        RECT 5.445 2.290 8.235 2.340 ;
        RECT 5.445 1.315 5.675 2.290 ;
        RECT 6.565 2.110 8.235 2.290 ;
        RECT 6.000 1.880 6.340 2.060 ;
        RECT 6.000 1.650 9.320 1.880 ;
        RECT 9.090 0.910 9.320 1.650 ;
        RECT 9.550 1.315 9.780 2.570 ;
        RECT 11.730 2.115 11.960 3.685 ;
        RECT 14.810 3.215 15.040 3.685 ;
        RECT 11.370 1.885 11.960 2.115 ;
        RECT 13.070 2.985 15.040 3.215 ;
        RECT 11.370 1.425 11.600 1.885 ;
        RECT 13.070 1.655 13.300 2.985 ;
        RECT 14.810 2.875 15.040 2.985 ;
        RECT 17.070 2.520 17.305 3.685 ;
        RECT 15.250 2.325 17.305 2.520 ;
        RECT 15.250 2.290 20.920 2.325 ;
        RECT 15.250 2.180 15.480 2.290 ;
        RECT 15.680 1.830 16.775 2.060 ;
        RECT 17.075 2.030 20.920 2.290 ;
        RECT 10.710 1.085 11.600 1.425 ;
        RECT 11.830 1.315 14.100 1.655 ;
        RECT 15.680 1.085 15.910 1.830 ;
        RECT 9.090 0.680 10.315 0.910 ;
        RECT 10.710 0.855 15.910 1.085 ;
        RECT 17.075 0.845 17.400 2.030 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffsnq_4
MACRO gf180mcu_fd_sc_mcu9t5v0__dlya_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlya_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.160 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 1.770 1.045 2.495 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.130 4.070 5.865 4.330 ;
        RECT 5.535 0.845 5.865 4.070 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 6.160 5.490 ;
        RECT 1.265 3.240 1.495 4.590 ;
        RECT 4.125 3.240 4.355 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.590 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.590 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.620 ;
        RECT 4.515 0.450 4.745 0.695 ;
        RECT 0.000 -0.450 6.160 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.955 0.475 3.580 ;
        RECT 0.245 2.725 2.035 2.955 ;
        RECT 0.245 1.280 0.475 2.725 ;
        RECT 1.805 1.740 2.035 2.725 ;
        RECT 2.385 2.495 2.615 3.580 ;
        RECT 3.105 3.010 3.335 3.580 ;
        RECT 3.105 2.780 4.290 3.010 ;
        RECT 4.060 2.585 4.290 2.780 ;
        RECT 2.385 1.795 3.830 2.495 ;
        RECT 2.385 1.280 2.715 1.795 ;
        RECT 4.060 1.745 5.185 2.585 ;
        RECT 4.055 1.695 5.185 1.745 ;
        RECT 4.055 0.910 4.285 1.695 ;
        RECT 3.000 0.680 4.285 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlya_1
MACRO gf180mcu_fd_sc_mcu9t5v0__dlya_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlya_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.210 0.970 2.795 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.130 3.265 5.615 4.330 ;
        RECT 5.130 3.035 6.435 3.265 ;
        RECT 6.205 1.990 6.435 3.035 ;
        RECT 5.485 1.760 6.435 1.990 ;
        RECT 5.485 0.845 5.715 1.760 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.280 5.490 ;
        RECT 1.265 3.485 1.495 4.590 ;
        RECT 4.130 3.485 4.360 4.590 ;
        RECT 6.505 3.485 6.735 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.645 ;
        RECT 4.365 0.450 4.595 0.960 ;
        RECT 6.625 0.450 6.855 1.630 ;
        RECT 0.000 -0.450 7.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.255 0.475 3.825 ;
        RECT 0.245 3.025 2.035 3.255 ;
        RECT 0.245 1.305 0.475 3.025 ;
        RECT 1.805 1.985 2.035 3.025 ;
        RECT 2.385 2.270 2.615 3.825 ;
        RECT 3.110 3.255 3.340 3.825 ;
        RECT 3.110 3.025 4.295 3.255 ;
        RECT 3.550 2.270 3.835 2.795 ;
        RECT 2.385 2.040 3.835 2.270 ;
        RECT 4.065 2.560 4.295 3.025 ;
        RECT 4.065 2.220 5.975 2.560 ;
        RECT 2.385 1.305 2.715 2.040 ;
        RECT 4.065 1.410 4.295 2.220 ;
        RECT 2.955 1.180 4.295 1.410 ;
        RECT 2.955 0.680 3.295 1.180 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlya_2
MACRO gf180mcu_fd_sc_mcu9t5v0__dlya_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlya_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.035 1.050 2.735 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.680 3.210 5.910 4.250 ;
        RECT 7.820 3.210 8.050 4.250 ;
        RECT 5.680 2.980 8.050 3.210 ;
        RECT 5.680 2.950 7.575 2.980 ;
        RECT 7.345 2.040 7.575 2.950 ;
        RECT 5.630 1.810 8.100 2.040 ;
        RECT 5.630 0.770 5.860 1.810 ;
        RECT 7.870 0.770 8.100 1.810 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 9.520 5.490 ;
        RECT 1.270 3.440 1.500 4.590 ;
        RECT 4.280 3.440 4.510 4.590 ;
        RECT 6.700 3.440 6.930 4.590 ;
        RECT 8.890 3.440 9.120 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.370 0.450 1.600 1.110 ;
        RECT 4.330 0.450 4.560 1.110 ;
        RECT 6.750 0.450 6.980 1.580 ;
        RECT 8.990 0.450 9.220 1.580 ;
        RECT 0.000 -0.450 9.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.250 3.195 0.480 3.780 ;
        RECT 0.250 2.965 2.095 3.195 ;
        RECT 0.250 0.770 0.480 2.965 ;
        RECT 1.755 2.035 2.095 2.965 ;
        RECT 2.390 2.735 2.620 3.780 ;
        RECT 3.260 3.210 3.490 3.780 ;
        RECT 3.260 2.980 4.445 3.210 ;
        RECT 2.390 2.505 3.985 2.735 ;
        RECT 3.700 2.030 3.985 2.505 ;
        RECT 2.490 1.800 3.985 2.030 ;
        RECT 4.215 2.500 4.445 2.980 ;
        RECT 4.215 2.270 7.115 2.500 ;
        RECT 2.490 0.770 2.720 1.800 ;
        RECT 4.215 1.570 4.445 2.270 ;
        RECT 3.210 1.340 4.445 1.570 ;
        RECT 3.210 0.770 3.440 1.340 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlya_4
MACRO gf180mcu_fd_sc_mcu9t5v0__dlyb_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyb_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 1.770 0.990 2.560 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.535 3.270 6.865 4.340 ;
        RECT 5.190 2.890 6.865 3.270 ;
        RECT 6.635 0.680 6.865 2.890 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.280 5.490 ;
        RECT 1.265 4.020 1.495 4.590 ;
        RECT 4.735 4.040 4.965 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.295 7.710 5.470 ;
        RECT -0.430 2.265 0.430 2.295 ;
        RECT 5.300 2.265 7.710 2.295 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 0.430 2.265 5.300 2.295 ;
        RECT -0.430 -0.430 7.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.965 ;
        RECT 4.835 0.450 5.065 0.695 ;
        RECT 0.000 -0.450 7.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 3.020 0.475 4.360 ;
        RECT 1.555 3.300 2.740 3.640 ;
        RECT 0.190 2.790 2.280 3.020 ;
        RECT 0.190 0.910 0.420 2.790 ;
        RECT 1.940 1.860 2.280 2.790 ;
        RECT 2.510 1.630 2.740 3.300 ;
        RECT 4.730 3.320 4.965 3.660 ;
        RECT 4.155 1.630 4.385 2.615 ;
        RECT 1.500 1.400 4.385 1.630 ;
        RECT 4.730 2.090 4.960 3.320 ;
        RECT 5.900 2.090 6.240 2.560 ;
        RECT 4.730 1.860 6.240 2.090 ;
        RECT 4.730 1.075 5.065 1.860 ;
        RECT 0.190 0.680 0.530 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyb_1
MACRO gf180mcu_fd_sc_mcu9t5v0__dlyb_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyb_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.400 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 1.770 0.990 2.560 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.912500 ;
    PORT
      LAYER Metal1 ;
        RECT 6.635 3.270 6.865 4.360 ;
        RECT 6.310 2.890 6.865 3.270 ;
        RECT 6.635 0.680 6.865 2.890 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 8.400 5.490 ;
        RECT 1.265 3.915 1.495 4.590 ;
        RECT 4.735 3.915 4.965 4.590 ;
        RECT 7.705 3.880 7.935 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.295 8.830 5.470 ;
        RECT -0.430 2.265 0.430 2.295 ;
        RECT 5.315 2.265 8.830 2.295 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 0.430 2.265 5.315 2.295 ;
        RECT -0.430 -0.430 8.830 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.965 ;
        RECT 4.835 0.450 5.065 0.695 ;
        RECT 7.755 0.450 7.985 1.435 ;
        RECT 0.000 -0.450 8.400 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 3.020 0.475 4.255 ;
        RECT 1.500 3.250 2.740 3.480 ;
        RECT 0.190 2.790 2.280 3.020 ;
        RECT 0.190 0.910 0.420 2.790 ;
        RECT 1.940 1.860 2.280 2.790 ;
        RECT 2.510 2.035 2.740 3.250 ;
        RECT 4.155 2.035 4.385 2.615 ;
        RECT 2.510 1.805 4.385 2.035 ;
        RECT 4.735 2.325 4.965 3.535 ;
        RECT 4.735 2.095 6.380 2.325 ;
        RECT 2.510 1.630 2.740 1.805 ;
        RECT 1.500 1.400 2.740 1.630 ;
        RECT 4.735 1.075 5.065 2.095 ;
        RECT 0.190 0.680 0.530 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyb_2
MACRO gf180mcu_fd_sc_mcu9t5v0__dlyb_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyb_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.640 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.900 0.970 2.710 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.825000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.740 3.650 6.970 4.360 ;
        RECT 8.930 3.650 9.160 4.360 ;
        RECT 6.740 3.420 9.160 3.650 ;
        RECT 8.930 1.590 9.160 3.420 ;
        RECT 6.690 1.210 9.160 1.590 ;
        RECT 6.690 0.680 6.920 1.210 ;
        RECT 8.930 0.680 9.160 1.210 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 10.640 5.490 ;
        RECT 1.320 4.060 1.550 4.590 ;
        RECT 4.790 4.060 5.020 4.590 ;
        RECT 7.760 3.880 7.990 4.590 ;
        RECT 9.950 3.880 10.180 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.295 11.070 5.470 ;
        RECT -0.430 2.265 0.430 2.295 ;
        RECT 5.370 2.265 11.070 2.295 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 0.430 2.265 5.370 2.295 ;
        RECT -0.430 -0.430 11.070 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.420 0.450 1.650 0.965 ;
        RECT 4.890 0.450 5.120 0.695 ;
        RECT 7.810 0.450 8.040 0.965 ;
        RECT 10.050 0.450 10.280 1.435 ;
        RECT 0.000 -0.450 10.640 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.170 0.585 4.345 ;
        RECT 1.555 3.395 2.795 3.625 ;
        RECT 0.245 2.940 1.505 3.170 ;
        RECT 0.245 0.910 0.475 2.940 ;
        RECT 1.275 2.655 1.505 2.940 ;
        RECT 1.275 2.425 2.335 2.655 ;
        RECT 2.050 1.900 2.335 2.425 ;
        RECT 2.565 1.630 2.795 3.395 ;
        RECT 4.210 1.630 4.440 2.710 ;
        RECT 1.555 1.400 4.440 1.630 ;
        RECT 4.790 2.420 5.020 3.680 ;
        RECT 4.790 2.190 8.175 2.420 ;
        RECT 4.790 1.075 5.120 2.190 ;
        RECT 0.245 0.680 0.585 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyb_4
MACRO gf180mcu_fd_sc_mcu9t5v0__dlyc_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyc_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.200 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 1.770 0.970 2.560 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.590 3.270 10.920 4.360 ;
        RECT 10.230 2.890 10.920 3.270 ;
        RECT 10.690 0.680 10.920 2.890 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 11.200 5.490 ;
        RECT 1.610 4.220 1.840 4.590 ;
        RECT 1.610 3.880 9.020 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.295 11.630 5.470 ;
        RECT -0.430 2.265 0.430 2.295 ;
        RECT 9.355 2.265 11.630 2.295 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 0.430 2.265 9.355 2.295 ;
        RECT -0.430 -0.430 11.630 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.965 ;
        RECT 4.890 0.450 5.120 0.690 ;
        RECT 8.890 0.450 9.120 0.695 ;
        RECT 0.000 -0.450 11.200 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.170 3.020 0.475 4.220 ;
        RECT 1.555 3.215 4.440 3.445 ;
        RECT 0.170 2.790 1.430 3.020 ;
        RECT 0.170 0.910 0.400 2.790 ;
        RECT 1.200 2.560 1.430 2.790 ;
        RECT 1.200 2.330 2.335 2.560 ;
        RECT 1.995 1.860 2.335 2.330 ;
        RECT 4.210 1.630 4.440 3.215 ;
        RECT 1.555 1.400 4.440 1.630 ;
        RECT 4.790 2.090 5.020 3.500 ;
        RECT 5.610 3.020 5.840 3.500 ;
        RECT 5.610 2.790 6.795 3.020 ;
        RECT 5.995 2.090 6.335 2.560 ;
        RECT 4.790 1.860 6.335 2.090 ;
        RECT 4.790 1.070 5.120 1.860 ;
        RECT 6.565 1.630 6.795 2.790 ;
        RECT 8.210 1.630 8.440 2.615 ;
        RECT 5.610 1.400 8.440 1.630 ;
        RECT 8.790 2.090 9.020 3.500 ;
        RECT 9.955 2.090 10.295 2.560 ;
        RECT 8.790 1.860 10.295 2.090 ;
        RECT 5.610 1.070 5.840 1.400 ;
        RECT 8.790 1.075 9.120 1.860 ;
        RECT 0.170 0.680 0.530 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyc_1
MACRO gf180mcu_fd_sc_mcu9t5v0__dlyc_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyc_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.320 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 1.770 0.990 2.560 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.912500 ;
    PORT
      LAYER Metal1 ;
        RECT 10.635 1.590 10.865 4.360 ;
        RECT 10.230 1.210 10.865 1.590 ;
        RECT 10.635 0.680 10.865 1.210 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 12.320 5.490 ;
        RECT 1.265 3.915 1.495 4.590 ;
        RECT 4.735 3.915 4.965 4.590 ;
        RECT 8.735 3.915 8.965 4.590 ;
        RECT 11.705 3.880 11.935 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.295 12.750 5.470 ;
        RECT -0.430 2.265 0.430 2.295 ;
        RECT 9.315 2.265 12.750 2.295 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 0.430 2.265 9.315 2.295 ;
        RECT -0.430 -0.430 12.750 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.965 ;
        RECT 4.835 0.450 5.065 0.690 ;
        RECT 8.835 0.450 9.065 0.695 ;
        RECT 11.755 0.450 11.985 1.435 ;
        RECT 0.000 -0.450 12.320 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 3.020 0.475 4.255 ;
        RECT 1.500 3.250 2.740 3.480 ;
        RECT 0.190 2.790 2.280 3.020 ;
        RECT 0.190 0.910 0.420 2.790 ;
        RECT 1.940 1.860 2.280 2.790 ;
        RECT 2.510 1.630 2.740 3.250 ;
        RECT 4.155 1.630 4.385 2.615 ;
        RECT 1.500 1.400 4.385 1.630 ;
        RECT 4.735 2.090 4.965 3.535 ;
        RECT 5.555 3.020 5.785 3.535 ;
        RECT 5.555 2.790 6.740 3.020 ;
        RECT 5.940 2.090 6.280 2.560 ;
        RECT 4.735 1.860 6.280 2.090 ;
        RECT 4.735 1.070 5.065 1.860 ;
        RECT 6.510 1.630 6.740 2.790 ;
        RECT 8.155 1.630 8.385 2.615 ;
        RECT 5.555 1.400 8.385 1.630 ;
        RECT 8.735 2.325 8.965 3.535 ;
        RECT 8.735 2.095 10.380 2.325 ;
        RECT 5.555 1.070 5.785 1.400 ;
        RECT 8.735 1.075 9.065 2.095 ;
        RECT 0.190 0.680 0.530 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyc_2
MACRO gf180mcu_fd_sc_mcu9t5v0__dlyc_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyc_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 1.140 0.990 1.840 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.565 3.105 10.795 3.685 ;
        RECT 12.705 3.105 12.935 3.685 ;
        RECT 10.565 2.875 12.935 3.105 ;
        RECT 12.225 1.655 12.455 2.875 ;
        RECT 10.565 1.425 13.035 1.655 ;
        RECT 10.565 0.845 10.795 1.425 ;
        RECT 12.470 0.845 13.035 1.425 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.560 5.490 ;
        RECT 1.265 3.710 1.495 4.590 ;
        RECT 4.665 3.710 4.895 4.590 ;
        RECT 8.665 3.710 8.895 4.590 ;
        RECT 11.585 3.875 11.815 4.590 ;
        RECT 13.825 3.875 14.055 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.380 14.990 5.470 ;
        RECT -0.430 2.265 0.430 2.380 ;
        RECT 9.065 2.265 14.990 2.380 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 0.430 2.265 9.065 2.380 ;
        RECT -0.430 -0.430 14.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.965 ;
        RECT 4.765 0.450 4.995 0.935 ;
        RECT 8.765 0.450 8.995 0.935 ;
        RECT 11.685 0.450 11.915 1.165 ;
        RECT 13.925 0.450 14.155 1.165 ;
        RECT 0.000 -0.450 14.560 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 2.760 0.475 4.050 ;
        RECT 1.485 2.990 4.315 3.330 ;
        RECT 0.190 2.530 2.210 2.760 ;
        RECT 0.190 0.910 0.420 2.530 ;
        RECT 1.870 2.060 2.210 2.530 ;
        RECT 4.085 1.715 4.315 2.990 ;
        RECT 1.430 1.485 4.315 1.715 ;
        RECT 4.665 2.060 4.895 3.330 ;
        RECT 5.485 2.990 5.715 3.330 ;
        RECT 5.485 2.760 8.315 2.990 ;
        RECT 5.870 2.060 6.210 2.530 ;
        RECT 4.665 1.830 6.210 2.060 ;
        RECT 4.665 1.315 4.995 1.830 ;
        RECT 8.085 1.600 8.315 2.760 ;
        RECT 5.430 1.370 8.315 1.600 ;
        RECT 8.665 2.315 8.895 3.330 ;
        RECT 8.665 1.975 11.995 2.315 ;
        RECT 8.665 1.315 8.995 1.975 ;
        RECT 0.190 0.680 0.530 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyc_4
MACRO gf180mcu_fd_sc_mcu9t5v0__dlyd_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyd_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.120 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 0.970 2.580 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.545 0.840 14.970 4.360 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 15.120 5.490 ;
        RECT 1.270 3.895 1.500 4.590 ;
        RECT 4.740 3.895 4.970 4.590 ;
        RECT 8.740 3.895 8.970 4.590 ;
        RECT 12.745 3.895 12.975 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.295 15.550 5.470 ;
        RECT -0.430 2.265 0.430 2.295 ;
        RECT 13.310 2.265 15.550 2.295 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 0.430 2.265 13.310 2.295 ;
        RECT -0.430 -0.430 15.550 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.370 0.450 1.600 0.965 ;
        RECT 4.840 0.450 5.070 0.930 ;
        RECT 8.840 0.450 9.070 0.930 ;
        RECT 12.845 0.450 13.075 0.690 ;
        RECT 0.000 -0.450 15.120 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.195 3.040 0.480 4.235 ;
        RECT 1.505 3.230 2.690 3.460 ;
        RECT 0.195 3.000 1.375 3.040 ;
        RECT 0.195 2.810 2.230 3.000 ;
        RECT 0.195 0.910 0.425 2.810 ;
        RECT 1.245 2.770 2.230 2.810 ;
        RECT 2.000 2.190 2.230 2.770 ;
        RECT 2.460 1.630 2.690 3.230 ;
        RECT 4.740 2.580 4.970 3.515 ;
        RECT 5.560 3.040 5.790 3.515 ;
        RECT 5.560 2.810 6.690 3.040 ;
        RECT 4.160 1.630 4.390 2.580 ;
        RECT 1.505 1.400 4.390 1.630 ;
        RECT 4.740 2.350 6.230 2.580 ;
        RECT 4.740 1.310 5.070 2.350 ;
        RECT 6.000 1.770 6.230 2.350 ;
        RECT 5.505 1.540 5.845 1.595 ;
        RECT 6.460 1.540 6.690 2.810 ;
        RECT 8.740 2.580 8.970 3.515 ;
        RECT 9.560 3.040 9.790 3.515 ;
        RECT 9.560 2.810 10.690 3.040 ;
        RECT 8.160 1.540 8.390 2.580 ;
        RECT 5.505 1.310 8.390 1.540 ;
        RECT 8.740 2.350 10.230 2.580 ;
        RECT 8.740 1.310 9.070 2.350 ;
        RECT 10.000 1.770 10.230 2.350 ;
        RECT 9.505 1.540 9.845 1.595 ;
        RECT 10.460 1.540 10.690 2.810 ;
        RECT 12.165 1.540 12.395 2.580 ;
        RECT 9.505 1.310 12.395 1.540 ;
        RECT 12.745 2.000 12.975 3.515 ;
        RECT 13.965 2.000 14.195 2.580 ;
        RECT 12.745 1.770 14.195 2.000 ;
        RECT 12.745 1.070 13.075 1.770 ;
        RECT 0.195 0.680 0.535 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyd_1
MACRO gf180mcu_fd_sc_mcu9t5v0__dlyd_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyd_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.240 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 1.770 0.990 2.570 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.530 4.070 14.765 4.360 ;
        RECT 14.535 3.365 14.765 4.070 ;
        RECT 14.535 3.135 15.585 3.365 ;
        RECT 15.355 1.820 15.585 3.135 ;
        RECT 14.635 1.590 15.585 1.820 ;
        RECT 14.635 0.845 14.865 1.590 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 16.240 5.490 ;
        RECT 1.265 3.925 1.495 4.590 ;
        RECT 4.735 3.925 4.965 4.590 ;
        RECT 8.735 3.925 8.965 4.590 ;
        RECT 12.735 3.925 12.965 4.590 ;
        RECT 15.655 3.585 15.885 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.295 16.670 5.470 ;
        RECT -0.430 2.265 0.430 2.295 ;
        RECT 13.315 2.265 16.670 2.295 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 0.430 2.265 13.315 2.295 ;
        RECT -0.430 -0.430 16.670 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.965 ;
        RECT 4.835 0.450 5.065 0.690 ;
        RECT 8.835 0.450 9.065 0.920 ;
        RECT 12.835 0.450 13.065 0.695 ;
        RECT 15.755 0.450 15.985 1.435 ;
        RECT 0.000 -0.450 16.240 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 3.030 0.475 4.265 ;
        RECT 1.500 3.260 4.385 3.490 ;
        RECT 0.190 2.800 2.225 3.030 ;
        RECT 0.190 0.910 0.420 2.800 ;
        RECT 1.995 2.220 2.225 2.800 ;
        RECT 4.155 1.630 4.385 3.260 ;
        RECT 1.500 1.400 4.385 1.630 ;
        RECT 4.735 2.625 4.965 3.545 ;
        RECT 5.555 3.085 5.785 3.545 ;
        RECT 5.555 2.855 8.385 3.085 ;
        RECT 4.735 1.815 6.225 2.625 ;
        RECT 4.735 1.070 5.065 1.815 ;
        RECT 8.155 1.585 8.385 2.855 ;
        RECT 5.555 1.355 8.385 1.585 ;
        RECT 8.735 2.625 8.965 3.545 ;
        RECT 9.555 3.085 9.785 3.545 ;
        RECT 9.555 2.855 12.385 3.085 ;
        RECT 8.735 1.815 10.225 2.625 ;
        RECT 5.555 1.070 5.785 1.355 ;
        RECT 8.735 1.300 9.065 1.815 ;
        RECT 12.155 1.585 12.385 2.855 ;
        RECT 9.500 1.355 12.385 1.585 ;
        RECT 12.735 2.390 12.965 3.545 ;
        RECT 12.735 2.050 15.125 2.390 ;
        RECT 12.735 1.075 13.065 2.050 ;
        RECT 0.190 0.680 0.530 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyd_2
MACRO gf180mcu_fd_sc_mcu9t5v0__dlyd_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyd_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.660 1.770 1.000 2.595 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.825000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.695 3.120 14.970 4.360 ;
        RECT 16.735 3.120 16.965 4.360 ;
        RECT 14.695 2.890 16.965 3.120 ;
        RECT 16.360 1.900 16.590 2.890 ;
        RECT 14.645 1.670 17.115 1.900 ;
        RECT 14.645 0.680 14.875 1.670 ;
        RECT 16.885 0.680 17.115 1.670 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 18.480 5.490 ;
        RECT 1.275 3.930 1.505 4.590 ;
        RECT 4.745 3.930 4.975 4.590 ;
        RECT 8.745 3.930 8.975 4.590 ;
        RECT 12.745 3.930 12.975 4.590 ;
        RECT 15.715 3.880 15.945 4.590 ;
        RECT 17.905 3.880 18.135 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.300 18.910 5.470 ;
        RECT -0.430 2.265 0.430 2.300 ;
        RECT 13.310 2.265 18.910 2.300 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 0.430 2.265 13.310 2.300 ;
        RECT -0.430 -0.430 18.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.375 0.450 1.605 0.970 ;
        RECT 4.845 0.450 5.075 0.970 ;
        RECT 8.845 0.450 9.075 0.965 ;
        RECT 12.845 0.450 13.075 0.695 ;
        RECT 15.765 0.450 15.995 1.440 ;
        RECT 18.005 0.450 18.235 1.440 ;
        RECT 0.000 -0.450 18.480 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.200 3.055 0.485 4.270 ;
        RECT 1.510 3.265 2.750 3.495 ;
        RECT 0.200 3.035 1.415 3.055 ;
        RECT 0.200 2.825 2.290 3.035 ;
        RECT 0.200 0.915 0.430 2.825 ;
        RECT 1.320 2.805 2.290 2.825 ;
        RECT 1.950 1.895 2.290 2.805 ;
        RECT 2.520 1.635 2.750 3.265 ;
        RECT 4.165 1.635 4.395 2.650 ;
        RECT 1.510 1.405 4.395 1.635 ;
        RECT 4.745 2.125 4.975 3.550 ;
        RECT 5.565 3.055 5.795 3.550 ;
        RECT 5.565 2.825 6.750 3.055 ;
        RECT 5.950 2.125 6.290 2.595 ;
        RECT 4.745 1.895 6.290 2.125 ;
        RECT 4.745 1.350 5.075 1.895 ;
        RECT 6.520 1.635 6.750 2.825 ;
        RECT 8.165 1.635 8.395 2.650 ;
        RECT 5.510 1.405 8.395 1.635 ;
        RECT 8.745 2.125 8.975 3.550 ;
        RECT 9.565 3.055 9.795 3.550 ;
        RECT 9.565 2.825 10.750 3.055 ;
        RECT 9.950 2.125 10.290 2.595 ;
        RECT 8.745 1.895 10.290 2.125 ;
        RECT 10.520 2.070 10.750 2.825 ;
        RECT 12.165 2.070 12.395 2.650 ;
        RECT 8.745 1.345 9.075 1.895 ;
        RECT 10.520 1.840 12.395 2.070 ;
        RECT 12.745 2.360 12.975 3.550 ;
        RECT 12.745 2.130 16.130 2.360 ;
        RECT 10.520 1.630 10.750 1.840 ;
        RECT 9.510 1.400 10.750 1.630 ;
        RECT 12.745 1.075 13.075 2.130 ;
        RECT 0.200 0.685 0.540 0.915 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyd_4
MACRO gf180mcu_fd_sc_mcu9t5v0__endcap
  CLASS ENDCAP PRE ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__endcap ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.120 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Nwell ;
        RECT -2.930 2.265 1.550 5.470 ;
      LAYER Metal1 ;
        RECT 0.000 4.590 1.120 5.490 ;
        RECT 0.230 2.340 0.850 4.590 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Pwell ;
        RECT -2.930 -0.430 1.550 2.265 ;
      LAYER Metal1 ;
        RECT 0.230 0.450 0.850 1.530 ;
        RECT 0.000 -0.450 1.120 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__endcap
MACRO gf180mcu_fd_sc_mcu9t5v0__fill_1
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fill_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 0.560 5.490 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 0.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 0.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.450 0.560 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__fill_1
MACRO gf180mcu_fd_sc_mcu9t5v0__fill_2
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fill_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.120 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 1.120 5.490 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 1.550 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 1.550 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.450 1.120 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__fill_2
MACRO gf180mcu_fd_sc_mcu9t5v0__fill_4
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fill_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 2.240 5.490 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 2.670 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.450 2.240 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__fill_4
MACRO gf180mcu_fd_sc_mcu9t5v0__fill_8
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fill_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 4.480 5.490 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.450 4.480 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__fill_8
MACRO gf180mcu_fd_sc_mcu9t5v0__fill_16
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fill_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.960 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 8.960 5.490 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.390 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.390 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.450 8.960 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__fill_16
MACRO gf180mcu_fd_sc_mcu9t5v0__fill_32
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fill_32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.920 5.490 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 18.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.450 17.920 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__fill_32
MACRO gf180mcu_fd_sc_mcu9t5v0__fill_64
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fill_64 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 35.840 5.490 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 36.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 36.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.450 35.840 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__fill_64
MACRO gf180mcu_fd_sc_mcu9t5v0__fillcap_4
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fillcap_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 2.240 5.490 ;
        RECT 1.765 3.550 1.995 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 2.670 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 0.000 -0.450 2.240 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.060 0.475 4.360 ;
        RECT 1.270 2.470 1.995 2.700 ;
        RECT 0.245 1.830 0.970 2.060 ;
        RECT 1.765 0.680 1.995 2.470 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__fillcap_4
MACRO gf180mcu_fd_sc_mcu9t5v0__fillcap_8
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fillcap_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 4.480 5.490 ;
        RECT 1.765 3.550 1.995 4.590 ;
        RECT 4.005 3.550 4.235 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 0.000 -0.450 4.480 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.060 0.475 4.360 ;
        RECT 1.270 2.470 1.995 2.700 ;
        RECT 0.245 1.830 0.970 2.060 ;
        RECT 1.765 0.680 1.995 2.470 ;
        RECT 2.485 2.060 2.715 4.360 ;
        RECT 3.510 2.470 4.235 2.700 ;
        RECT 2.485 1.830 3.210 2.060 ;
        RECT 4.005 0.680 4.235 2.470 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__fillcap_8
MACRO gf180mcu_fd_sc_mcu9t5v0__fillcap_16
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fillcap_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.960 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 8.960 5.490 ;
        RECT 1.765 3.550 1.995 4.590 ;
        RECT 4.005 3.550 4.235 4.590 ;
        RECT 6.245 3.550 6.475 4.590 ;
        RECT 8.485 3.550 8.715 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.390 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.390 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 6.965 0.450 7.195 1.490 ;
        RECT 0.000 -0.450 8.960 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.060 0.475 4.360 ;
        RECT 1.270 2.470 1.995 2.700 ;
        RECT 0.245 1.830 0.970 2.060 ;
        RECT 1.765 0.680 1.995 2.470 ;
        RECT 2.485 2.060 2.715 4.360 ;
        RECT 3.510 2.470 4.235 2.700 ;
        RECT 2.485 1.830 3.210 2.060 ;
        RECT 4.005 0.680 4.235 2.470 ;
        RECT 4.725 2.060 4.955 4.360 ;
        RECT 5.750 2.470 6.475 2.700 ;
        RECT 4.725 1.830 5.450 2.060 ;
        RECT 6.245 0.680 6.475 2.470 ;
        RECT 6.965 2.060 7.195 4.360 ;
        RECT 7.990 2.470 8.715 2.700 ;
        RECT 6.965 1.830 7.690 2.060 ;
        RECT 8.485 0.680 8.715 2.470 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__fillcap_16
MACRO gf180mcu_fd_sc_mcu9t5v0__fillcap_32
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fillcap_32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.920 5.490 ;
        RECT 1.765 3.550 1.995 4.590 ;
        RECT 4.005 3.550 4.235 4.590 ;
        RECT 6.245 3.550 6.475 4.590 ;
        RECT 8.485 3.550 8.715 4.590 ;
        RECT 10.725 3.550 10.955 4.590 ;
        RECT 12.965 3.550 13.195 4.590 ;
        RECT 15.205 3.550 15.435 4.590 ;
        RECT 17.445 3.550 17.675 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 18.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 6.965 0.450 7.195 1.490 ;
        RECT 9.205 0.450 9.435 1.490 ;
        RECT 11.445 0.450 11.675 1.490 ;
        RECT 13.685 0.450 13.915 1.490 ;
        RECT 15.925 0.450 16.155 1.490 ;
        RECT 0.000 -0.450 17.920 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.060 0.475 4.360 ;
        RECT 0.245 1.830 0.970 2.060 ;
        RECT 1.325 1.490 1.555 2.755 ;
        RECT 2.485 2.060 2.715 4.360 ;
        RECT 2.485 1.830 3.210 2.060 ;
        RECT 3.565 1.490 3.795 2.755 ;
        RECT 4.725 2.060 4.955 4.360 ;
        RECT 4.725 1.830 5.450 2.060 ;
        RECT 5.805 1.490 6.035 2.755 ;
        RECT 6.965 2.060 7.195 4.360 ;
        RECT 6.965 1.830 7.690 2.060 ;
        RECT 8.045 1.490 8.275 2.755 ;
        RECT 9.205 2.060 9.435 4.360 ;
        RECT 9.205 1.830 9.930 2.060 ;
        RECT 10.285 1.490 10.515 2.755 ;
        RECT 11.445 2.060 11.675 4.360 ;
        RECT 11.445 1.830 12.170 2.060 ;
        RECT 12.525 1.490 12.755 2.755 ;
        RECT 13.685 2.060 13.915 4.360 ;
        RECT 13.685 1.830 14.410 2.060 ;
        RECT 14.765 1.490 14.995 2.755 ;
        RECT 15.925 2.060 16.155 4.360 ;
        RECT 15.925 1.830 16.650 2.060 ;
        RECT 17.005 1.490 17.235 2.755 ;
        RECT 1.325 1.260 1.995 1.490 ;
        RECT 3.565 1.260 4.235 1.490 ;
        RECT 5.805 1.260 6.475 1.490 ;
        RECT 8.045 1.260 8.715 1.490 ;
        RECT 10.285 1.260 10.955 1.490 ;
        RECT 12.525 1.260 13.195 1.490 ;
        RECT 14.765 1.260 15.435 1.490 ;
        RECT 17.005 1.260 17.675 1.490 ;
        RECT 1.765 0.680 1.995 1.260 ;
        RECT 4.005 0.680 4.235 1.260 ;
        RECT 6.245 0.680 6.475 1.260 ;
        RECT 8.485 0.680 8.715 1.260 ;
        RECT 10.725 0.680 10.955 1.260 ;
        RECT 12.965 0.680 13.195 1.260 ;
        RECT 15.205 0.680 15.435 1.260 ;
        RECT 17.445 0.680 17.675 1.260 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__fillcap_32
MACRO gf180mcu_fd_sc_mcu9t5v0__fillcap_64
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fillcap_64 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 35.840 5.490 ;
        RECT 1.765 3.550 1.995 4.590 ;
        RECT 4.005 3.550 4.235 4.590 ;
        RECT 6.245 3.550 6.475 4.590 ;
        RECT 8.485 3.550 8.715 4.590 ;
        RECT 10.725 3.550 10.955 4.590 ;
        RECT 12.965 3.550 13.195 4.590 ;
        RECT 15.205 3.550 15.435 4.590 ;
        RECT 17.445 3.550 17.675 4.590 ;
        RECT 19.685 3.550 19.915 4.590 ;
        RECT 21.925 3.550 22.155 4.590 ;
        RECT 24.165 3.550 24.395 4.590 ;
        RECT 26.405 3.550 26.635 4.590 ;
        RECT 28.645 3.550 28.875 4.590 ;
        RECT 30.885 3.550 31.115 4.590 ;
        RECT 33.125 3.550 33.355 4.590 ;
        RECT 35.365 3.550 35.595 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 36.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 36.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 6.965 0.450 7.195 1.490 ;
        RECT 9.205 0.450 9.435 1.490 ;
        RECT 11.445 0.450 11.675 1.490 ;
        RECT 13.685 0.450 13.915 1.490 ;
        RECT 15.925 0.450 16.155 1.490 ;
        RECT 18.165 0.450 18.395 1.490 ;
        RECT 20.405 0.450 20.635 1.490 ;
        RECT 22.645 0.450 22.875 1.490 ;
        RECT 24.885 0.450 25.115 1.490 ;
        RECT 27.125 0.450 27.355 1.490 ;
        RECT 29.365 0.450 29.595 1.490 ;
        RECT 31.605 0.450 31.835 1.490 ;
        RECT 33.845 0.450 34.075 1.490 ;
        RECT 0.000 -0.450 35.840 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.060 0.475 4.360 ;
        RECT 0.245 1.830 0.970 2.060 ;
        RECT 1.325 1.490 1.555 2.755 ;
        RECT 2.485 2.060 2.715 4.360 ;
        RECT 2.485 1.830 3.210 2.060 ;
        RECT 3.565 1.490 3.795 2.755 ;
        RECT 4.725 2.060 4.955 4.360 ;
        RECT 4.725 1.830 5.450 2.060 ;
        RECT 5.805 1.490 6.035 2.755 ;
        RECT 6.965 2.060 7.195 4.360 ;
        RECT 6.965 1.830 7.690 2.060 ;
        RECT 8.045 1.490 8.275 2.755 ;
        RECT 9.205 2.060 9.435 4.360 ;
        RECT 9.205 1.830 9.930 2.060 ;
        RECT 10.285 1.490 10.515 2.755 ;
        RECT 11.445 2.060 11.675 4.360 ;
        RECT 11.445 1.830 12.170 2.060 ;
        RECT 12.525 1.490 12.755 2.755 ;
        RECT 13.685 2.060 13.915 4.360 ;
        RECT 13.685 1.830 14.410 2.060 ;
        RECT 14.765 1.490 14.995 2.755 ;
        RECT 15.925 2.060 16.155 4.360 ;
        RECT 15.925 1.830 16.650 2.060 ;
        RECT 17.005 1.490 17.235 2.755 ;
        RECT 18.165 2.060 18.395 4.360 ;
        RECT 18.165 1.830 18.890 2.060 ;
        RECT 19.245 1.490 19.475 2.755 ;
        RECT 20.405 2.060 20.635 4.360 ;
        RECT 20.405 1.830 21.130 2.060 ;
        RECT 21.485 1.490 21.715 2.755 ;
        RECT 22.645 2.060 22.875 4.360 ;
        RECT 22.645 1.830 23.370 2.060 ;
        RECT 23.725 1.490 23.955 2.755 ;
        RECT 24.885 2.060 25.115 4.360 ;
        RECT 24.885 1.830 25.610 2.060 ;
        RECT 25.965 1.490 26.195 2.755 ;
        RECT 27.125 2.060 27.355 4.360 ;
        RECT 27.125 1.830 27.850 2.060 ;
        RECT 28.205 1.490 28.435 2.755 ;
        RECT 29.365 2.060 29.595 4.360 ;
        RECT 29.365 1.830 30.090 2.060 ;
        RECT 30.445 1.490 30.675 2.755 ;
        RECT 31.605 2.060 31.835 4.360 ;
        RECT 31.605 1.830 32.330 2.060 ;
        RECT 32.685 1.490 32.915 2.755 ;
        RECT 33.845 2.060 34.075 4.360 ;
        RECT 33.845 1.830 34.570 2.060 ;
        RECT 34.925 1.490 35.155 2.755 ;
        RECT 1.325 1.260 1.995 1.490 ;
        RECT 3.565 1.260 4.235 1.490 ;
        RECT 5.805 1.260 6.475 1.490 ;
        RECT 8.045 1.260 8.715 1.490 ;
        RECT 10.285 1.260 10.955 1.490 ;
        RECT 12.525 1.260 13.195 1.490 ;
        RECT 14.765 1.260 15.435 1.490 ;
        RECT 17.005 1.260 17.675 1.490 ;
        RECT 19.245 1.260 19.915 1.490 ;
        RECT 21.485 1.260 22.155 1.490 ;
        RECT 23.725 1.260 24.395 1.490 ;
        RECT 25.965 1.260 26.635 1.490 ;
        RECT 28.205 1.260 28.875 1.490 ;
        RECT 30.445 1.260 31.115 1.490 ;
        RECT 32.685 1.260 33.355 1.490 ;
        RECT 34.925 1.260 35.595 1.490 ;
        RECT 1.765 0.680 1.995 1.260 ;
        RECT 4.005 0.680 4.235 1.260 ;
        RECT 6.245 0.680 6.475 1.260 ;
        RECT 8.485 0.680 8.715 1.260 ;
        RECT 10.725 0.680 10.955 1.260 ;
        RECT 12.965 0.680 13.195 1.260 ;
        RECT 15.205 0.680 15.435 1.260 ;
        RECT 17.445 0.680 17.675 1.260 ;
        RECT 19.685 0.680 19.915 1.260 ;
        RECT 21.925 0.680 22.155 1.260 ;
        RECT 24.165 0.680 24.395 1.260 ;
        RECT 26.405 0.680 26.635 1.260 ;
        RECT 28.645 0.680 28.875 1.260 ;
        RECT 30.885 0.680 31.115 1.260 ;
        RECT 33.125 0.680 33.355 1.260 ;
        RECT 35.365 0.680 35.595 1.260 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__fillcap_64
MACRO gf180mcu_fd_sc_mcu9t5v0__filltie
  CLASS core WELLTAP ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__filltie ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.120 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 1.550 5.470 ;
      LAYER Metal1 ;
        RECT 0.000 4.590 1.120 5.490 ;
        RECT 0.330 2.340 0.710 4.590 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 1.550 2.265 ;
      LAYER Metal1 ;
        RECT 0.330 0.450 0.710 1.910 ;
        RECT 0.000 -0.450 1.120 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__filltie
MACRO gf180mcu_fd_sc_mcu9t5v0__hold
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__hold ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN Z
    DIRECTION INOUT ;
    ANTENNAGATEAREA 1.707000 ;
    ANTENNADIFFAREA 0.489600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 1.645 0.575 3.605 ;
        RECT 3.510 1.645 3.950 2.575 ;
        RECT 0.245 1.415 3.950 1.645 ;
        RECT 0.245 0.845 0.475 1.415 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.040 5.490 ;
        RECT 3.225 3.265 3.455 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 5.470 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 5.470 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.225 0.450 3.455 1.185 ;
        RECT 0.000 -0.450 5.040 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 4.245 3.035 4.575 4.075 ;
        RECT 2.510 2.805 4.575 3.035 ;
        RECT 2.510 1.875 2.850 2.805 ;
        RECT 4.345 0.845 4.575 2.805 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__hold
MACRO gf180mcu_fd_sc_mcu9t5v0__icgtn_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.800 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.350 1.770 11.715 2.710 ;
    END
  END CLKN
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.210 1.770 2.090 2.265 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.265 0.410 2.710 ;
        RECT 0.150 1.770 0.915 2.265 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.245200 ;
    PORT
      LAYER Metal1 ;
        RECT 16.195 3.830 16.475 4.200 ;
        RECT 15.830 3.390 16.475 3.830 ;
        RECT 16.245 1.590 16.475 3.390 ;
        RECT 15.830 1.210 16.475 1.590 ;
        RECT 16.245 0.795 16.475 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 16.800 5.490 ;
        RECT 0.675 3.390 0.905 4.590 ;
        RECT 5.805 3.390 6.035 4.590 ;
        RECT 8.665 3.390 8.895 4.590 ;
        RECT 12.245 3.390 12.475 4.590 ;
        RECT 15.175 3.390 15.405 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 17.230 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 17.230 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.080 ;
        RECT 5.805 0.450 6.035 1.135 ;
        RECT 8.765 0.450 8.995 1.135 ;
        RECT 12.165 0.450 12.395 1.135 ;
        RECT 14.405 0.450 14.635 1.135 ;
        RECT 15.125 0.450 15.355 1.605 ;
        RECT 0.000 -0.450 16.800 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.555 3.160 3.785 4.200 ;
        RECT 6.265 4.130 8.335 4.360 ;
        RECT 6.265 3.160 6.495 4.130 ;
        RECT 2.985 2.930 6.495 3.160 ;
        RECT 0.245 1.310 2.715 1.540 ;
        RECT 0.245 0.795 0.475 1.310 ;
        RECT 2.485 0.795 2.715 1.310 ;
        RECT 2.985 1.080 3.215 2.930 ;
        RECT 6.825 2.700 7.155 3.900 ;
        RECT 3.445 2.470 7.155 2.700 ;
        RECT 3.445 1.790 3.675 2.470 ;
        RECT 2.985 0.850 3.890 1.080 ;
        RECT 6.925 0.795 7.155 2.470 ;
        RECT 7.645 1.695 7.875 3.900 ;
        RECT 8.105 1.925 8.335 4.130 ;
        RECT 9.685 4.130 12.015 4.360 ;
        RECT 8.565 1.980 9.390 2.210 ;
        RECT 8.565 1.695 8.795 1.980 ;
        RECT 7.645 1.465 8.795 1.695 ;
        RECT 7.645 0.795 7.875 1.465 ;
        RECT 9.685 0.795 10.115 4.130 ;
        RECT 11.225 3.170 11.455 3.900 ;
        RECT 10.385 2.940 11.455 3.170 ;
        RECT 11.785 3.160 12.015 4.130 ;
        RECT 10.385 1.080 10.615 2.940 ;
        RECT 11.785 2.930 12.915 3.160 ;
        RECT 12.685 1.925 12.915 2.930 ;
        RECT 14.005 2.210 14.235 4.200 ;
        RECT 14.005 1.980 15.740 2.210 ;
        RECT 14.005 1.520 14.235 1.980 ;
        RECT 13.285 1.290 14.235 1.520 ;
        RECT 10.385 0.850 11.330 1.080 ;
        RECT 13.285 0.795 13.515 1.290 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtn_1
MACRO gf180mcu_fd_sc_mcu9t5v0__icgtn_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.640000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.350 1.770 11.675 2.710 ;
    END
  END CLKN
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.390 1.770 2.650 2.710 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 0.970 2.710 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.471600 ;
    PORT
      LAYER Metal1 ;
        RECT 16.275 0.815 16.650 4.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.920 5.490 ;
        RECT 1.435 3.400 1.665 4.590 ;
        RECT 5.805 3.400 6.035 4.590 ;
        RECT 8.625 3.400 8.855 4.590 ;
        RECT 12.025 3.400 12.255 4.590 ;
        RECT 15.255 3.400 15.485 4.590 ;
        RECT 17.295 3.400 17.525 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 18.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.100 ;
        RECT 5.565 0.450 5.795 1.155 ;
        RECT 8.525 0.450 8.755 1.155 ;
        RECT 11.925 0.450 12.155 1.155 ;
        RECT 14.165 0.450 14.395 1.155 ;
        RECT 15.205 0.450 15.435 1.625 ;
        RECT 17.445 0.450 17.675 1.625 ;
        RECT 0.000 -0.450 17.920 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 4.045 3.170 4.275 4.210 ;
        RECT 6.265 4.130 8.345 4.360 ;
        RECT 6.265 3.170 6.495 4.130 ;
        RECT 4.045 3.065 6.495 3.170 ;
        RECT 2.930 2.940 6.495 3.065 ;
        RECT 2.930 2.835 4.240 2.940 ;
        RECT 2.930 1.615 3.160 2.835 ;
        RECT 4.435 2.075 4.775 2.710 ;
        RECT 6.825 2.075 7.055 3.900 ;
        RECT 3.390 1.845 7.055 2.075 ;
        RECT 1.065 1.540 2.295 1.560 ;
        RECT 0.245 1.330 2.295 1.540 ;
        RECT 2.930 1.385 3.835 1.615 ;
        RECT 0.245 1.310 1.160 1.330 ;
        RECT 0.245 0.815 0.475 1.310 ;
        RECT 2.065 1.155 2.295 1.330 ;
        RECT 2.065 0.815 2.715 1.155 ;
        RECT 3.605 0.815 3.835 1.385 ;
        RECT 6.685 0.815 7.055 1.845 ;
        RECT 7.405 1.655 7.835 3.900 ;
        RECT 8.115 1.885 8.345 4.130 ;
        RECT 9.645 3.980 11.795 4.210 ;
        RECT 8.575 1.940 9.350 2.170 ;
        RECT 8.575 1.655 8.805 1.940 ;
        RECT 7.405 1.425 8.805 1.655 ;
        RECT 7.405 0.815 7.635 1.425 ;
        RECT 9.645 0.815 9.875 3.980 ;
        RECT 11.005 3.140 11.235 3.720 ;
        RECT 10.305 2.910 11.235 3.140 ;
        RECT 11.565 3.170 11.795 3.980 ;
        RECT 11.565 2.940 12.695 3.170 ;
        RECT 10.305 1.540 10.535 2.910 ;
        RECT 12.465 2.415 12.695 2.940 ;
        RECT 13.785 2.170 14.015 4.210 ;
        RECT 13.785 1.940 15.980 2.170 ;
        RECT 13.785 1.560 14.015 1.940 ;
        RECT 10.305 1.310 11.090 1.540 ;
        RECT 12.990 1.330 14.015 1.560 ;
        RECT 12.990 1.310 13.330 1.330 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtn_2
MACRO gf180mcu_fd_sc_mcu9t5v0__icgtn_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtn_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.160 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.640000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.350 1.770 11.610 2.710 ;
    END
  END CLKN
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.345 1.820 2.650 3.270 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 0.970 2.710 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.943200 ;
    PORT
      LAYER Metal1 ;
        RECT 16.030 2.920 16.260 3.960 ;
        RECT 18.070 2.920 18.550 3.960 ;
        RECT 16.030 2.690 18.550 2.920 ;
        RECT 18.070 1.600 18.550 2.690 ;
        RECT 16.030 1.300 18.550 1.600 ;
        RECT 16.030 0.790 16.310 1.300 ;
        RECT 18.320 0.790 18.550 1.300 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 20.160 5.490 ;
        RECT 1.325 3.150 1.555 4.590 ;
        RECT 5.820 3.150 6.050 4.590 ;
        RECT 8.580 3.150 8.810 4.590 ;
        RECT 12.080 3.785 12.310 4.590 ;
        RECT 15.010 3.150 15.240 4.590 ;
        RECT 17.050 3.150 17.280 4.590 ;
        RECT 19.090 3.150 19.320 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 20.590 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 20.590 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.075 ;
        RECT 5.580 0.450 5.810 1.130 ;
        RECT 8.580 0.450 8.810 1.130 ;
        RECT 11.980 0.450 12.210 1.130 ;
        RECT 14.220 0.450 14.450 1.130 ;
        RECT 14.960 0.450 15.190 1.600 ;
        RECT 17.200 0.450 17.430 1.070 ;
        RECT 19.440 0.450 19.670 1.600 ;
        RECT 0.000 -0.450 20.160 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 6.280 4.130 8.250 4.360 ;
        RECT 4.060 2.920 4.290 3.960 ;
        RECT 6.280 2.920 6.510 4.130 ;
        RECT 4.060 2.795 6.510 2.920 ;
        RECT 2.945 2.690 6.510 2.795 ;
        RECT 2.945 2.565 4.265 2.690 ;
        RECT 2.945 1.615 3.175 2.565 ;
        RECT 4.470 2.075 4.810 2.460 ;
        RECT 6.840 2.075 7.070 3.900 ;
        RECT 3.405 1.845 7.070 2.075 ;
        RECT 0.245 1.305 2.715 1.535 ;
        RECT 2.945 1.385 3.850 1.615 ;
        RECT 0.245 0.790 0.475 1.305 ;
        RECT 2.485 0.790 2.715 1.305 ;
        RECT 3.620 0.790 3.850 1.385 ;
        RECT 6.700 0.790 7.070 1.845 ;
        RECT 7.460 1.590 7.790 3.900 ;
        RECT 8.020 1.820 8.250 4.130 ;
        RECT 9.600 3.735 9.830 3.960 ;
        RECT 9.600 3.555 11.855 3.735 ;
        RECT 9.600 3.505 12.750 3.555 ;
        RECT 8.480 1.875 9.305 2.105 ;
        RECT 8.480 1.590 8.710 1.875 ;
        RECT 7.460 1.360 8.710 1.590 ;
        RECT 7.460 0.790 7.690 1.360 ;
        RECT 9.600 0.790 9.930 3.505 ;
        RECT 11.630 3.325 12.750 3.505 ;
        RECT 10.860 2.935 11.290 3.275 ;
        RECT 10.360 1.460 10.590 2.200 ;
        RECT 10.860 1.460 11.090 2.935 ;
        RECT 12.520 2.475 12.750 3.325 ;
        RECT 13.840 2.320 14.070 3.960 ;
        RECT 13.840 1.980 17.510 2.320 ;
        RECT 13.840 1.535 14.070 1.980 ;
        RECT 10.360 1.230 11.090 1.460 ;
        RECT 13.045 1.305 14.070 1.535 ;
        RECT 13.045 1.285 13.385 1.305 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtn_4
MACRO gf180mcu_fd_sc_mcu9t5v0__icgtp_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.120 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.230 1.770 10.490 2.710 ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.255 2.710 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.270 1.190 2.500 ;
        RECT 0.150 1.210 0.410 2.270 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.245200 ;
    PORT
      LAYER Metal1 ;
        RECT 14.150 0.695 14.610 3.685 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 15.120 5.490 ;
        RECT 0.845 3.435 1.075 4.590 ;
        RECT 6.025 3.910 6.255 4.590 ;
        RECT 8.980 4.235 9.210 4.590 ;
        RECT 8.980 4.005 13.240 4.235 ;
        RECT 8.980 3.895 11.200 4.005 ;
        RECT 13.010 3.425 13.240 4.005 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 15.550 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 15.550 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.530 0.450 1.870 1.075 ;
        RECT 5.785 0.450 6.015 1.130 ;
        RECT 9.260 0.450 9.490 1.035 ;
        RECT 13.260 0.450 13.490 1.015 ;
        RECT 0.000 -0.450 15.120 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.205 3.175 3.595 4.245 ;
        RECT 7.045 3.640 7.275 4.245 ;
        RECT 5.680 3.410 10.975 3.640 ;
        RECT 3.205 2.945 5.450 3.175 ;
        RECT 0.640 1.305 2.935 1.535 ;
        RECT 0.640 0.980 0.870 1.305 ;
        RECT 0.190 0.750 0.870 0.980 ;
        RECT 2.705 0.790 2.935 1.305 ;
        RECT 3.205 1.075 3.435 2.945 ;
        RECT 3.665 2.485 4.990 2.715 ;
        RECT 3.665 1.790 3.895 2.485 ;
        RECT 5.220 1.985 5.450 2.945 ;
        RECT 5.680 2.215 5.910 3.410 ;
        RECT 6.140 2.270 6.750 2.500 ;
        RECT 6.140 1.985 6.370 2.270 ;
        RECT 5.220 1.755 6.370 1.985 ;
        RECT 6.980 1.130 7.210 3.410 ;
        RECT 8.135 2.605 8.475 3.180 ;
        RECT 7.565 2.375 8.475 2.605 ;
        RECT 9.770 2.950 10.515 3.180 ;
        RECT 9.770 2.500 10.000 2.950 ;
        RECT 3.205 0.845 4.110 1.075 ;
        RECT 6.905 0.790 7.210 1.130 ;
        RECT 8.140 0.695 8.475 2.375 ;
        RECT 8.715 2.270 10.000 2.500 ;
        RECT 10.745 2.500 10.975 3.410 ;
        RECT 11.990 3.105 12.220 3.685 ;
        RECT 11.990 2.875 13.015 3.105 ;
        RECT 12.785 2.500 13.015 2.875 ;
        RECT 10.745 2.270 12.555 2.500 ;
        RECT 12.785 2.270 13.915 2.500 ;
        RECT 9.770 0.980 10.000 2.270 ;
        RECT 12.785 1.035 13.015 2.270 ;
        RECT 9.770 0.750 10.665 0.980 ;
        RECT 11.100 0.695 13.015 1.035 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtp_1
MACRO gf180mcu_fd_sc_mcu9t5v0__icgtp_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.680 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.625000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.230 1.210 10.490 2.405 ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.210 1.770 2.090 2.350 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 0.970 2.710 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.471600 ;
    PORT
      LAYER Metal1 ;
        RECT 13.590 2.890 14.200 3.685 ;
        RECT 13.940 1.590 14.200 2.890 ;
        RECT 13.590 1.210 14.200 1.590 ;
        RECT 13.940 0.790 14.200 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 15.680 5.490 ;
        RECT 0.695 3.440 0.925 4.590 ;
        RECT 5.805 3.850 6.035 4.590 ;
        RECT 8.720 4.250 8.950 4.590 ;
        RECT 8.720 4.020 15.220 4.250 ;
        RECT 8.720 3.850 11.140 4.020 ;
        RECT 12.950 3.440 13.180 4.020 ;
        RECT 14.990 3.440 15.220 4.020 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 16.110 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 16.110 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.075 ;
        RECT 5.620 0.450 5.850 1.130 ;
        RECT 9.020 0.450 9.250 1.130 ;
        RECT 12.820 0.450 13.050 1.430 ;
        RECT 15.060 0.450 15.290 1.430 ;
        RECT 0.000 -0.450 15.680 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.555 3.175 3.785 4.250 ;
        RECT 6.825 3.620 7.055 4.250 ;
        RECT 5.460 3.390 11.700 3.620 ;
        RECT 2.985 2.945 5.230 3.175 ;
        RECT 0.245 1.305 2.715 1.535 ;
        RECT 0.245 0.790 0.475 1.305 ;
        RECT 2.485 0.790 2.715 1.305 ;
        RECT 2.985 1.075 3.215 2.945 ;
        RECT 3.445 2.485 4.770 2.715 ;
        RECT 3.445 1.790 3.675 2.485 ;
        RECT 5.000 1.835 5.230 2.945 ;
        RECT 5.460 2.065 5.690 3.390 ;
        RECT 6.005 1.835 6.345 2.350 ;
        RECT 5.000 1.605 6.345 1.835 ;
        RECT 2.985 0.845 3.890 1.075 ;
        RECT 6.740 0.790 6.970 3.390 ;
        RECT 7.400 2.930 7.985 3.160 ;
        RECT 9.685 2.930 10.025 3.160 ;
        RECT 7.400 1.075 7.630 2.930 ;
        RECT 9.685 2.350 9.915 2.930 ;
        RECT 8.225 2.120 9.915 2.350 ;
        RECT 11.470 2.350 11.700 3.390 ;
        RECT 11.930 3.105 12.160 3.685 ;
        RECT 11.930 2.875 12.885 3.105 ;
        RECT 12.655 2.405 12.885 2.875 ;
        RECT 11.470 2.120 12.425 2.350 ;
        RECT 7.400 0.845 8.185 1.075 ;
        RECT 9.685 0.980 9.915 2.120 ;
        RECT 12.655 2.065 13.490 2.405 ;
        RECT 12.655 1.890 12.885 2.065 ;
        RECT 10.860 1.660 12.885 1.890 ;
        RECT 9.685 0.750 10.425 0.980 ;
        RECT 10.860 0.790 11.090 1.660 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtp_2
MACRO gf180mcu_fd_sc_mcu9t5v0__icgtp_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.625000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.230 1.770 10.490 2.710 ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.405 0.970 2.710 ;
        RECT 0.710 2.175 2.090 2.405 ;
        RECT 0.710 1.770 0.970 2.175 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.110000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 1.770 0.415 2.710 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.943200 ;
    PORT
      LAYER Metal1 ;
        RECT 13.885 3.105 14.145 3.685 ;
        RECT 15.955 3.105 16.355 3.685 ;
        RECT 13.885 2.875 16.355 3.105 ;
        RECT 15.955 1.745 16.355 2.875 ;
        RECT 13.885 1.515 16.355 1.745 ;
        RECT 13.885 0.795 14.115 1.515 ;
        RECT 15.770 0.710 16.355 1.515 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.920 5.490 ;
        RECT 0.625 3.440 0.855 4.590 ;
        RECT 5.805 3.855 6.035 4.590 ;
        RECT 8.865 3.855 9.095 4.590 ;
        RECT 10.855 3.855 11.085 4.590 ;
        RECT 12.895 4.250 13.125 4.590 ;
        RECT 12.895 4.020 17.205 4.250 ;
        RECT 12.895 3.440 13.125 4.020 ;
        RECT 14.935 3.440 15.165 4.020 ;
        RECT 16.975 3.440 17.205 4.020 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 18.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.080 ;
        RECT 5.565 0.450 5.795 1.135 ;
        RECT 8.965 0.450 9.195 1.135 ;
        RECT 12.765 0.450 12.995 1.485 ;
        RECT 15.005 0.450 15.235 1.035 ;
        RECT 17.245 0.450 17.475 1.485 ;
        RECT 0.000 -0.450 17.920 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 4.035 3.230 4.265 4.250 ;
        RECT 6.825 3.625 7.055 4.250 ;
        RECT 5.405 3.395 11.645 3.625 ;
        RECT 4.035 3.050 5.175 3.230 ;
        RECT 2.985 3.000 5.175 3.050 ;
        RECT 2.985 2.820 4.260 3.000 ;
        RECT 0.245 1.310 2.715 1.540 ;
        RECT 0.245 0.795 0.475 1.310 ;
        RECT 2.485 0.795 2.715 1.310 ;
        RECT 2.985 1.080 3.215 2.820 ;
        RECT 4.485 2.130 4.715 2.770 ;
        RECT 3.445 1.790 4.715 2.130 ;
        RECT 4.945 1.890 5.175 3.000 ;
        RECT 5.405 2.120 5.635 3.395 ;
        RECT 5.865 2.175 6.530 2.405 ;
        RECT 5.865 1.890 6.095 2.175 ;
        RECT 4.945 1.660 6.095 1.890 ;
        RECT 6.760 1.135 6.990 3.395 ;
        RECT 7.790 2.460 8.130 3.160 ;
        RECT 7.345 2.120 8.130 2.460 ;
        RECT 9.770 2.935 10.170 3.165 ;
        RECT 9.770 2.405 10.000 2.935 ;
        RECT 8.370 2.175 10.000 2.405 ;
        RECT 11.415 2.405 11.645 3.395 ;
        RECT 11.875 3.105 12.105 3.685 ;
        RECT 11.875 2.875 13.060 3.105 ;
        RECT 11.415 2.175 12.600 2.405 ;
        RECT 12.830 2.315 13.060 2.875 ;
        RECT 2.985 0.850 3.890 1.080 ;
        RECT 6.685 0.795 6.990 1.135 ;
        RECT 7.845 0.795 8.130 2.120 ;
        RECT 9.770 1.540 10.000 2.175 ;
        RECT 12.830 1.975 15.370 2.315 ;
        RECT 12.830 1.945 13.060 1.975 ;
        RECT 10.805 1.715 13.060 1.945 ;
        RECT 9.770 1.310 10.315 1.540 ;
        RECT 10.085 0.795 10.315 1.310 ;
        RECT 10.805 0.795 11.035 1.715 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtp_4
MACRO gf180mcu_fd_sc_mcu9t5v0__inv_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.300 1.070 2.530 ;
        RECT 0.710 1.210 1.015 2.300 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 2.150 1.595 4.360 ;
        RECT 1.270 0.680 1.595 2.150 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 2.240 5.490 ;
        RECT 0.345 3.550 0.575 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 2.670 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 0.000 -0.450 2.240 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_1
MACRO gf180mcu_fd_sc_mcu9t5v0__inv_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 2.270 1.910 2.710 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.915500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.395 3.830 1.625 4.360 ;
        RECT 1.395 3.450 2.370 3.830 ;
        RECT 2.140 1.850 2.370 3.450 ;
        RECT 1.830 1.670 2.370 1.850 ;
        RECT 1.830 1.490 2.285 1.670 ;
        RECT 1.395 1.210 2.285 1.490 ;
        RECT 1.395 0.680 1.625 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 3.360 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.600 3.550 2.830 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 3.790 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 3.790 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.515 0.450 2.745 1.490 ;
        RECT 0.000 -0.450 3.360 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_2
MACRO gf180mcu_fd_sc_mcu9t5v0__inv_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.121000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.410 2.270 2.160 2.710 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.207000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 1.365 3.090 3.735 3.320 ;
        RECT 2.390 1.950 2.805 3.090 ;
        RECT 1.365 1.720 3.835 1.950 ;
        RECT 1.365 0.680 1.595 1.720 ;
        RECT 3.605 0.680 3.835 1.720 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 4.480 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 0.000 -0.450 4.480 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_3
MACRO gf180mcu_fd_sc_mcu9t5v0__inv_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.580 2.270 2.330 2.650 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.350 1.595 4.360 ;
        RECT 3.505 3.350 3.835 4.360 ;
        RECT 1.365 3.120 3.835 3.350 ;
        RECT 3.335 1.890 3.835 3.120 ;
        RECT 1.365 1.660 3.835 1.890 ;
        RECT 1.365 0.680 1.595 1.660 ;
        RECT 3.605 0.680 3.835 1.660 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.600 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.580 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.430 ;
        RECT 2.485 0.450 2.715 1.430 ;
        RECT 4.725 0.450 4.955 1.430 ;
        RECT 0.000 -0.450 5.600 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_4
MACRO gf180mcu_fd_sc_mcu9t5v0__inv_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 13.655999 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 2.265 4.260 2.645 ;
        RECT 5.360 2.215 8.880 2.650 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.284000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 5.745 3.320 5.975 4.360 ;
        RECT 7.985 3.320 8.215 4.360 ;
        RECT 1.365 3.090 8.215 3.320 ;
        RECT 4.630 1.985 5.130 3.090 ;
        RECT 1.365 1.755 8.315 1.985 ;
        RECT 1.365 0.680 1.595 1.755 ;
        RECT 3.575 0.680 3.835 1.755 ;
        RECT 5.845 0.680 6.075 1.755 ;
        RECT 8.085 0.680 8.315 1.755 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 10.080 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 10.510 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.165 ;
        RECT 6.965 0.450 7.195 1.490 ;
        RECT 9.205 0.450 9.435 1.490 ;
        RECT 0.000 -0.450 10.080 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_8
MACRO gf180mcu_fd_sc_mcu9t5v0__inv_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 20.483999 ;
    PORT
      LAYER Metal1 ;
        RECT 0.180 2.270 5.690 2.650 ;
        RECT 7.600 2.215 13.000 2.650 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 10.926000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 5.745 3.320 5.975 4.360 ;
        RECT 7.985 3.320 8.215 4.360 ;
        RECT 10.225 3.320 10.455 4.360 ;
        RECT 12.465 3.320 12.695 4.360 ;
        RECT 1.365 3.090 12.695 3.320 ;
        RECT 6.755 1.950 7.370 3.090 ;
        RECT 1.365 1.720 12.795 1.950 ;
        RECT 1.365 0.680 1.625 1.720 ;
        RECT 3.605 0.680 3.835 1.720 ;
        RECT 5.845 0.680 6.075 1.720 ;
        RECT 8.085 0.680 8.315 1.720 ;
        RECT 10.325 0.680 10.555 1.720 ;
        RECT 12.565 0.680 12.795 1.720 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.560 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
        RECT 11.345 3.550 11.575 4.590 ;
        RECT 13.585 3.550 13.815 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 6.965 0.450 7.195 1.490 ;
        RECT 9.205 0.450 9.435 1.490 ;
        RECT 11.445 0.450 11.675 1.490 ;
        RECT 13.685 0.450 13.915 1.490 ;
        RECT 0.000 -0.450 14.560 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_12
MACRO gf180mcu_fd_sc_mcu9t5v0__inv_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 27.311998 ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 2.215 7.965 2.650 ;
        RECT 9.225 2.215 16.505 2.650 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 14.568000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.210 1.595 4.360 ;
        RECT 3.505 3.210 3.735 4.360 ;
        RECT 5.745 3.210 5.975 4.360 ;
        RECT 8.080 3.210 8.310 4.360 ;
        RECT 1.365 3.180 8.310 3.210 ;
        RECT 10.225 3.180 10.455 4.360 ;
        RECT 12.465 3.180 12.695 4.360 ;
        RECT 14.705 3.180 14.935 4.360 ;
        RECT 16.945 3.180 17.175 4.360 ;
        RECT 1.365 2.980 17.175 3.180 ;
        RECT 8.195 2.950 17.175 2.980 ;
        RECT 8.195 1.950 8.995 2.950 ;
        RECT 1.365 1.720 17.275 1.950 ;
        RECT 1.365 0.680 1.625 1.720 ;
        RECT 3.605 0.680 3.835 1.720 ;
        RECT 5.845 0.680 6.075 1.720 ;
        RECT 8.085 0.680 8.315 1.720 ;
        RECT 10.325 0.680 10.555 1.720 ;
        RECT 12.565 0.680 12.795 1.720 ;
        RECT 14.805 0.680 15.035 1.720 ;
        RECT 17.045 0.680 17.275 1.720 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 19.040 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
        RECT 11.345 3.550 11.575 4.590 ;
        RECT 13.585 3.550 13.815 4.590 ;
        RECT 15.825 3.550 16.055 4.590 ;
        RECT 18.065 3.550 18.295 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 19.470 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 19.470 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 6.965 0.450 7.195 1.490 ;
        RECT 9.205 0.450 9.435 1.490 ;
        RECT 11.445 0.450 11.675 1.490 ;
        RECT 13.685 0.450 13.915 1.490 ;
        RECT 15.925 0.450 16.155 1.490 ;
        RECT 18.165 0.450 18.395 1.490 ;
        RECT 0.000 -0.450 19.040 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_16
MACRO gf180mcu_fd_sc_mcu9t5v0__inv_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_20 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 34.139999 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 2.270 9.900 2.650 ;
        RECT 11.110 2.270 20.380 2.650 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 18.209999 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.320 1.595 4.360 ;
        RECT 3.505 3.320 3.735 4.360 ;
        RECT 5.745 3.320 5.975 4.360 ;
        RECT 7.985 3.320 8.215 4.360 ;
        RECT 10.225 3.320 10.455 4.360 ;
        RECT 12.465 3.320 12.695 4.360 ;
        RECT 14.705 3.320 14.935 4.360 ;
        RECT 16.945 3.320 17.175 4.360 ;
        RECT 19.185 3.320 19.415 4.360 ;
        RECT 21.425 3.320 21.655 4.360 ;
        RECT 1.365 3.090 21.655 3.320 ;
        RECT 10.130 1.950 10.880 3.090 ;
        RECT 1.335 1.720 21.755 1.950 ;
        RECT 1.335 0.680 1.595 1.720 ;
        RECT 3.605 0.680 3.835 1.720 ;
        RECT 5.845 0.680 6.075 1.720 ;
        RECT 8.085 0.680 8.315 1.720 ;
        RECT 10.325 0.680 10.555 1.720 ;
        RECT 12.565 0.680 12.795 1.720 ;
        RECT 14.805 0.680 15.035 1.720 ;
        RECT 17.045 0.680 17.275 1.720 ;
        RECT 19.285 0.680 19.515 1.720 ;
        RECT 21.525 0.680 21.755 1.720 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 23.520 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
        RECT 9.105 3.550 9.335 4.590 ;
        RECT 11.345 3.550 11.575 4.590 ;
        RECT 13.585 3.550 13.815 4.590 ;
        RECT 15.825 3.550 16.055 4.590 ;
        RECT 18.065 3.550 18.295 4.590 ;
        RECT 20.305 3.550 20.535 4.590 ;
        RECT 22.545 3.550 22.775 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 23.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 23.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 6.965 0.450 7.195 1.490 ;
        RECT 9.205 0.450 9.435 1.490 ;
        RECT 11.445 0.450 11.675 1.490 ;
        RECT 13.685 0.450 13.915 1.490 ;
        RECT 15.925 0.450 16.155 1.490 ;
        RECT 18.165 0.450 18.395 1.490 ;
        RECT 20.405 0.450 20.635 1.490 ;
        RECT 22.645 0.450 22.875 1.490 ;
        RECT 0.000 -0.450 23.520 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_20
MACRO gf180mcu_fd_sc_mcu9t5v0__invz_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.698000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.015 0.970 2.710 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.849000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.505 1.770 8.810 2.710 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.372800 ;
    PORT
      LAYER Metal1 ;
        RECT 4.610 1.770 4.890 3.900 ;
        RECT 4.610 1.140 4.840 1.770 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 9.520 5.490 ;
        RECT 1.265 3.480 1.495 4.590 ;
        RECT 5.680 3.860 5.910 4.590 ;
        RECT 7.585 3.480 7.815 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.610 0.450 1.840 1.480 ;
        RECT 5.730 0.450 5.960 1.165 ;
        RECT 7.585 0.450 7.815 1.480 ;
        RECT 0.000 -0.450 9.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.250 0.475 4.290 ;
        RECT 2.335 4.130 5.350 4.360 ;
        RECT 2.335 3.480 2.565 4.130 ;
        RECT 0.245 3.020 3.060 3.250 ;
        RECT 2.105 2.245 2.335 3.020 ;
        RECT 1.200 2.015 2.335 2.245 ;
        RECT 1.200 1.820 1.430 2.015 ;
        RECT 1.095 1.625 1.430 1.820 ;
        RECT 1.095 1.425 1.325 1.625 ;
        RECT 3.355 1.425 3.585 3.820 ;
        RECT 0.190 1.195 1.325 1.425 ;
        RECT 2.675 1.195 3.585 1.425 ;
        RECT 3.355 0.910 3.585 1.195 ;
        RECT 3.850 1.140 4.080 4.130 ;
        RECT 5.120 3.630 5.350 4.130 ;
        RECT 6.565 3.630 6.795 4.290 ;
        RECT 5.120 3.400 6.795 3.630 ;
        RECT 5.120 2.430 5.415 3.400 ;
        RECT 8.945 3.380 9.175 4.290 ;
        RECT 8.045 3.150 9.175 3.380 ;
        RECT 8.045 2.245 8.275 3.150 ;
        RECT 5.145 1.625 5.375 2.170 ;
        RECT 7.090 2.015 8.275 2.245 ;
        RECT 5.145 1.565 6.695 1.625 ;
        RECT 5.070 1.395 6.695 1.565 ;
        RECT 5.070 0.910 5.300 1.395 ;
        RECT 6.465 1.140 6.695 1.395 ;
        RECT 8.045 1.425 8.275 2.015 ;
        RECT 8.045 1.195 9.330 1.425 ;
        RECT 3.355 0.680 5.300 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_1
MACRO gf180mcu_fd_sc_mcu9t5v0__invz_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 0.970 2.710 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.692000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.990 1.770 8.460 2.710 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.622400 ;
    PORT
      LAYER Metal1 ;
        RECT 6.770 2.710 7.000 3.750 ;
        RECT 6.770 1.490 7.130 2.710 ;
        RECT 6.620 1.210 7.130 1.490 ;
        RECT 6.620 0.680 6.850 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 9.520 5.490 ;
        RECT 1.370 3.400 1.600 4.590 ;
        RECT 5.750 4.350 5.980 4.590 ;
        RECT 7.790 3.400 8.020 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.420 0.450 1.650 1.020 ;
        RECT 5.500 0.450 5.730 1.020 ;
        RECT 7.740 0.450 7.970 1.490 ;
        RECT 0.000 -0.450 9.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.350 3.170 0.580 4.210 ;
        RECT 2.900 4.130 4.960 4.360 ;
        RECT 2.900 3.400 3.130 4.130 ;
        RECT 0.350 2.940 3.625 3.170 ;
        RECT 1.860 2.470 3.625 2.940 ;
        RECT 1.860 1.490 2.090 2.470 ;
        RECT 3.920 2.240 4.150 3.900 ;
        RECT 3.200 2.010 4.150 2.240 ;
        RECT 4.585 2.220 4.960 4.130 ;
        RECT 6.165 3.980 7.560 4.210 ;
        RECT 6.165 3.155 6.395 3.980 ;
        RECT 5.240 2.925 6.395 3.155 ;
        RECT 7.330 3.170 7.560 3.980 ;
        RECT 8.810 3.170 9.090 4.210 ;
        RECT 7.330 2.940 9.090 3.170 ;
        RECT 5.240 2.450 5.470 2.925 ;
        RECT 5.700 2.465 6.475 2.695 ;
        RECT 5.700 2.220 5.930 2.465 ;
        RECT 3.200 1.490 3.430 2.010 ;
        RECT 4.585 1.990 5.930 2.220 ;
        RECT 4.585 1.780 4.815 1.990 ;
        RECT 0.300 1.260 2.090 1.490 ;
        RECT 0.300 0.680 0.530 1.260 ;
        RECT 2.540 1.085 3.430 1.490 ;
        RECT 3.660 1.550 4.815 1.780 ;
        RECT 3.660 1.315 3.890 1.550 ;
        RECT 6.160 1.480 6.390 2.110 ;
        RECT 5.035 1.250 6.390 1.480 ;
        RECT 5.035 1.085 5.265 1.250 ;
        RECT 2.540 0.680 5.265 1.085 ;
        RECT 8.860 0.680 9.090 2.940 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_2
MACRO gf180mcu_fd_sc_mcu9t5v0__invz_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.880 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 0.970 2.710 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.692000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.190 1.770 5.645 2.710 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.995200 ;
    PORT
      LAYER Metal1 ;
        RECT 9.465 3.195 9.930 4.210 ;
        RECT 11.505 3.195 11.735 4.210 ;
        RECT 9.465 2.965 12.495 3.195 ;
        RECT 12.265 1.600 12.495 2.965 ;
        RECT 10.025 1.370 12.495 1.600 ;
        RECT 10.025 0.790 10.255 1.370 ;
        RECT 12.265 0.840 12.495 1.370 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 12.880 5.490 ;
        RECT 1.370 3.845 1.600 4.590 ;
        RECT 6.045 4.280 6.275 4.590 ;
        RECT 8.265 3.400 8.495 4.590 ;
        RECT 10.485 3.880 10.715 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 13.310 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.310 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.420 0.450 1.650 1.020 ;
        RECT 6.235 0.450 6.575 0.620 ;
        RECT 8.725 0.450 8.955 1.160 ;
        RECT 11.145 0.450 11.375 1.020 ;
        RECT 0.000 -0.450 12.880 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.350 3.170 0.580 4.210 ;
        RECT 2.895 4.050 5.825 4.210 ;
        RECT 2.895 3.980 7.475 4.050 ;
        RECT 2.895 3.400 3.125 3.980 ;
        RECT 0.350 2.940 3.565 3.170 ;
        RECT 3.335 2.060 3.565 2.940 ;
        RECT 1.200 1.830 3.565 2.060 ;
        RECT 3.795 2.940 4.145 3.750 ;
        RECT 1.200 1.540 1.430 1.830 ;
        RECT 0.300 1.310 1.430 1.540 ;
        RECT 3.795 1.490 4.025 2.940 ;
        RECT 4.375 1.655 4.605 3.980 ;
        RECT 5.605 3.820 7.475 3.980 ;
        RECT 5.025 3.170 5.255 3.750 ;
        RECT 5.025 2.940 6.980 3.170 ;
        RECT 0.300 0.680 0.530 1.310 ;
        RECT 2.540 1.080 4.025 1.490 ;
        RECT 4.255 1.315 4.605 1.655 ;
        RECT 6.750 2.060 6.980 2.940 ;
        RECT 7.245 2.735 7.475 3.820 ;
        RECT 7.245 2.505 11.365 2.735 ;
        RECT 6.750 1.540 7.090 2.060 ;
        RECT 4.920 1.310 7.090 1.540 ;
        RECT 7.605 1.830 12.030 2.060 ;
        RECT 7.605 1.080 7.835 1.830 ;
        RECT 2.540 0.850 7.835 1.080 ;
        RECT 2.540 0.680 2.770 0.850 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_3
MACRO gf180mcu_fd_sc_mcu9t5v0__invz_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.440 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.060 0.410 2.710 ;
        RECT 0.150 1.770 1.020 2.060 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.692000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.130 1.830 6.070 2.650 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.244800 ;
    PORT
      LAYER Metal1 ;
        RECT 9.110 3.310 9.410 3.900 ;
        RECT 11.190 3.310 11.870 3.900 ;
        RECT 9.110 2.965 11.870 3.310 ;
        RECT 11.585 1.620 11.870 2.965 ;
        RECT 9.180 1.390 11.870 1.620 ;
        RECT 9.180 0.730 9.630 1.390 ;
        RECT 11.640 0.730 11.870 1.390 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 13.440 5.490 ;
        RECT 1.315 3.845 1.545 4.590 ;
        RECT 6.040 3.800 6.270 4.590 ;
        RECT 8.130 3.880 8.360 4.590 ;
        RECT 10.170 3.880 10.400 4.590 ;
        RECT 12.210 3.090 12.440 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 13.870 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.870 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.070 ;
        RECT 5.985 0.450 6.325 0.635 ;
        RECT 8.280 0.450 8.510 0.690 ;
        RECT 10.520 0.450 10.750 1.160 ;
        RECT 12.760 0.450 12.990 1.540 ;
        RECT 0.000 -0.450 13.440 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.925 4.130 5.810 4.360 ;
        RECT 0.295 3.320 0.525 3.900 ;
        RECT 0.295 3.090 1.480 3.320 ;
        RECT 2.925 3.090 3.155 4.130 ;
        RECT 1.250 2.060 1.480 3.090 ;
        RECT 3.365 2.520 3.595 2.755 ;
        RECT 1.860 2.290 3.595 2.520 ;
        RECT 1.860 2.060 2.090 2.290 ;
        RECT 3.945 2.060 4.175 3.900 ;
        RECT 1.250 1.830 2.090 2.060 ;
        RECT 3.090 1.830 4.175 2.060 ;
        RECT 1.250 1.540 1.480 1.830 ;
        RECT 0.245 1.310 1.480 1.540 ;
        RECT 0.245 0.730 0.475 1.310 ;
        RECT 2.485 0.960 2.715 1.540 ;
        RECT 3.090 1.135 3.320 1.830 ;
        RECT 4.405 1.600 4.635 4.130 ;
        RECT 5.020 3.110 5.250 3.900 ;
        RECT 5.580 3.570 5.810 4.130 ;
        RECT 7.110 3.570 7.345 4.150 ;
        RECT 5.580 3.340 7.345 3.570 ;
        RECT 5.020 2.880 6.760 3.110 ;
        RECT 3.550 1.370 4.635 1.600 ;
        RECT 6.530 1.595 6.760 2.880 ;
        RECT 7.115 2.735 7.345 3.340 ;
        RECT 7.115 2.505 11.075 2.735 ;
        RECT 4.865 1.365 6.760 1.595 ;
        RECT 8.720 1.850 10.265 2.110 ;
        RECT 8.720 1.270 8.950 1.850 ;
        RECT 7.235 1.135 8.950 1.270 ;
        RECT 3.090 1.040 8.950 1.135 ;
        RECT 3.090 0.960 7.445 1.040 ;
        RECT 2.485 0.905 7.445 0.960 ;
        RECT 2.485 0.730 3.315 0.905 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_4
MACRO gf180mcu_fd_sc_mcu9t5v0__invz_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.720 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 1.770 1.555 2.710 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.165 2.330 5.450 3.270 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.669600 ;
    PORT
      LAYER Metal1 ;
        RECT 12.215 3.155 12.455 4.190 ;
        RECT 14.255 3.155 14.485 4.190 ;
        RECT 16.295 3.155 16.525 4.195 ;
        RECT 18.335 3.155 18.805 4.195 ;
        RECT 12.215 2.925 18.805 3.155 ;
        RECT 18.315 1.595 18.805 2.925 ;
        RECT 12.165 1.215 19.115 1.595 ;
        RECT 12.165 1.210 14.635 1.215 ;
        RECT 12.165 0.680 12.395 1.210 ;
        RECT 14.405 0.680 14.635 1.210 ;
        RECT 16.645 1.210 19.115 1.215 ;
        RECT 16.645 0.680 16.875 1.210 ;
        RECT 18.885 0.680 19.115 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 20.720 5.490 ;
        RECT 1.905 3.420 2.135 4.590 ;
        RECT 4.675 4.350 4.905 4.590 ;
        RECT 6.715 4.350 6.945 4.590 ;
        RECT 8.755 3.380 8.985 4.590 ;
        RECT 10.995 3.880 11.225 4.590 ;
        RECT 13.235 3.385 13.465 4.590 ;
        RECT 15.275 3.385 15.505 4.590 ;
        RECT 17.315 3.385 17.545 4.590 ;
        RECT 19.355 3.380 19.585 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 21.150 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.150 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.020 ;
        RECT 4.270 0.450 4.610 0.635 ;
        RECT 6.510 0.450 6.850 0.635 ;
        RECT 8.805 0.450 9.035 1.490 ;
        RECT 11.045 0.450 11.275 1.490 ;
        RECT 13.285 0.450 13.515 0.980 ;
        RECT 15.525 0.450 15.755 0.980 ;
        RECT 17.765 0.450 17.995 0.980 ;
        RECT 20.005 0.450 20.235 1.490 ;
        RECT 0.000 -0.450 20.720 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.885 3.170 1.115 4.190 ;
        RECT 7.735 4.120 7.965 4.190 ;
        RECT 2.925 3.890 7.965 4.120 ;
        RECT 2.925 3.380 3.155 3.890 ;
        RECT 0.885 3.150 2.725 3.170 ;
        RECT 0.885 2.940 3.650 3.150 ;
        RECT 2.630 2.425 3.650 2.940 ;
        RECT 2.630 2.110 2.860 2.425 ;
        RECT 1.805 1.880 2.860 2.110 ;
        RECT 3.945 2.055 4.175 3.660 ;
        RECT 1.805 1.490 2.035 1.880 ;
        RECT 3.090 1.825 4.175 2.055 ;
        RECT 3.090 1.490 3.320 1.825 ;
        RECT 4.405 1.595 4.635 3.890 ;
        RECT 5.695 2.710 5.925 3.660 ;
        RECT 5.695 2.480 7.385 2.710 ;
        RECT 7.155 1.595 7.385 2.480 ;
        RECT 7.735 2.695 7.965 3.890 ;
        RECT 9.875 2.695 10.105 4.190 ;
        RECT 7.735 2.405 17.195 2.695 ;
        RECT 0.245 1.260 2.035 1.490 ;
        RECT 0.245 0.680 0.475 1.260 ;
        RECT 2.485 1.135 3.320 1.490 ;
        RECT 3.550 1.365 4.635 1.595 ;
        RECT 5.390 1.365 7.385 1.595 ;
        RECT 7.745 1.825 17.535 2.055 ;
        RECT 7.745 1.135 7.975 1.825 ;
        RECT 2.485 0.905 7.975 1.135 ;
        RECT 2.485 0.680 2.715 0.905 ;
        RECT 7.630 0.855 7.975 0.905 ;
        RECT 9.925 0.840 10.155 1.825 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_8
MACRO gf180mcu_fd_sc_mcu9t5v0__invz_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 29.120 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 0.970 2.710 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.076000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.570 1.785 6.010 3.270 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 10.274400 ;
    PORT
      LAYER Metal1 ;
        RECT 16.140 3.490 16.370 4.280 ;
        RECT 18.280 3.490 18.510 4.280 ;
        RECT 20.520 3.490 20.750 4.280 ;
        RECT 22.660 3.490 22.890 4.280 ;
        RECT 24.700 3.490 24.930 4.280 ;
        RECT 26.735 3.490 26.970 4.280 ;
        RECT 16.140 3.010 26.970 3.490 ;
        RECT 26.450 1.595 26.980 3.010 ;
        RECT 16.090 0.895 27.520 1.595 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 29.120 5.490 ;
        RECT 1.830 3.470 2.060 4.590 ;
        RECT 6.030 4.510 6.260 4.590 ;
        RECT 8.510 4.510 8.740 4.590 ;
        RECT 10.770 3.950 11.000 4.590 ;
        RECT 12.810 3.470 13.040 4.590 ;
        RECT 14.920 3.880 15.150 4.590 ;
        RECT 17.160 3.960 17.390 4.590 ;
        RECT 19.400 3.940 19.630 4.590 ;
        RECT 21.640 3.940 21.870 4.590 ;
        RECT 23.680 3.940 23.910 4.590 ;
        RECT 25.720 3.940 25.950 4.590 ;
        RECT 27.760 3.470 27.990 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 29.550 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 29.550 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.070 ;
        RECT 5.955 0.450 6.295 0.635 ;
        RECT 8.195 0.450 8.535 0.635 ;
        RECT 10.490 0.450 10.720 1.540 ;
        RECT 12.730 0.450 12.960 1.540 ;
        RECT 14.970 0.450 15.200 1.540 ;
        RECT 17.155 0.450 17.495 0.635 ;
        RECT 19.395 0.450 19.735 0.635 ;
        RECT 21.635 0.450 21.975 0.635 ;
        RECT 23.875 0.450 24.215 0.635 ;
        RECT 26.115 0.450 26.455 0.635 ;
        RECT 28.410 0.450 28.640 1.540 ;
        RECT 0.000 -0.450 29.120 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.810 3.170 1.040 4.280 ;
        RECT 2.850 4.050 9.980 4.280 ;
        RECT 2.850 3.470 3.080 4.050 ;
        RECT 0.810 2.940 3.575 3.170 ;
        RECT 1.805 2.480 3.575 2.940 ;
        RECT 1.805 1.540 2.035 2.480 ;
        RECT 3.870 2.055 4.100 3.820 ;
        RECT 3.090 1.825 4.100 2.055 ;
        RECT 0.245 1.310 2.035 1.540 ;
        RECT 0.245 0.730 0.475 1.310 ;
        RECT 2.485 1.095 2.715 1.540 ;
        RECT 3.090 1.095 3.320 1.825 ;
        RECT 4.330 1.595 4.560 4.050 ;
        RECT 4.790 3.590 7.500 3.820 ;
        RECT 4.790 3.010 5.020 3.590 ;
        RECT 7.270 2.525 7.500 3.590 ;
        RECT 9.750 2.735 9.980 4.050 ;
        RECT 11.790 2.735 12.020 4.280 ;
        RECT 13.830 2.735 14.060 4.280 ;
        RECT 7.270 2.230 8.975 2.525 ;
        RECT 9.750 2.505 25.570 2.735 ;
        RECT 3.550 1.365 4.560 1.595 ;
        RECT 8.690 1.555 8.975 2.230 ;
        RECT 4.835 1.325 8.975 1.555 ;
        RECT 9.430 1.825 25.940 2.055 ;
        RECT 9.430 1.095 9.660 1.825 ;
        RECT 2.485 0.865 9.660 1.095 ;
        RECT 2.485 0.730 2.715 0.865 ;
        RECT 9.315 0.815 9.660 0.865 ;
        RECT 11.610 0.840 11.840 1.825 ;
        RECT 13.850 0.840 14.080 1.825 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_12
MACRO gf180mcu_fd_sc_mcu9t5v0__invz_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 36.960 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.815 1.850 1.155 2.275 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.768000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.065 2.030 7.710 2.605 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 14.329200 ;
    PORT
      LAYER Metal1 ;
        RECT 19.405 3.365 19.635 4.120 ;
        RECT 21.545 3.365 21.775 4.120 ;
        RECT 23.785 3.365 24.015 4.120 ;
        RECT 26.025 3.365 26.255 4.120 ;
        RECT 28.265 3.365 28.495 4.120 ;
        RECT 30.505 3.365 30.735 4.120 ;
        RECT 32.745 3.365 32.975 4.120 ;
        RECT 35.085 3.365 35.315 4.120 ;
        RECT 19.405 2.965 35.315 3.365 ;
        RECT 34.835 1.595 35.315 2.965 ;
        RECT 19.405 0.895 35.315 1.595 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 36.960 5.490 ;
        RECT 1.905 3.310 2.135 4.590 ;
        RECT 4.665 4.350 4.895 4.590 ;
        RECT 6.805 4.350 7.035 4.590 ;
        RECT 9.045 3.310 9.275 4.590 ;
        RECT 11.285 3.310 11.515 4.590 ;
        RECT 13.525 3.310 13.755 4.590 ;
        RECT 15.765 3.310 15.995 4.590 ;
        RECT 18.185 3.880 18.415 4.590 ;
        RECT 20.425 3.745 20.655 4.590 ;
        RECT 22.665 3.745 22.895 4.590 ;
        RECT 24.905 3.745 25.135 4.590 ;
        RECT 27.145 3.745 27.375 4.590 ;
        RECT 29.385 3.745 29.615 4.590 ;
        RECT 31.625 3.745 31.855 4.590 ;
        RECT 33.865 3.745 34.095 4.590 ;
        RECT 36.105 3.310 36.335 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 37.390 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 37.390 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.160 ;
        RECT 4.610 0.450 4.950 0.640 ;
        RECT 6.850 0.450 7.190 0.640 ;
        RECT 9.090 0.450 9.430 0.640 ;
        RECT 11.385 0.450 11.615 1.455 ;
        RECT 13.625 0.450 13.855 1.490 ;
        RECT 15.865 0.450 16.095 1.490 ;
        RECT 18.285 0.450 18.515 1.490 ;
        RECT 20.470 0.450 20.810 0.665 ;
        RECT 22.710 0.450 23.050 0.665 ;
        RECT 24.950 0.450 25.290 0.665 ;
        RECT 27.190 0.450 27.530 0.665 ;
        RECT 29.430 0.450 29.770 0.665 ;
        RECT 31.670 0.450 32.010 0.665 ;
        RECT 33.910 0.450 34.250 0.665 ;
        RECT 36.205 0.450 36.435 1.490 ;
        RECT 0.000 -0.450 36.960 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.885 2.735 1.115 4.120 ;
        RECT 2.925 3.890 8.815 4.120 ;
        RECT 2.925 3.310 3.155 3.890 ;
        RECT 0.885 2.505 3.650 2.735 ;
        RECT 1.805 1.620 2.035 2.505 ;
        RECT 3.945 2.095 4.175 3.650 ;
        RECT 0.245 1.390 2.035 1.620 ;
        RECT 3.090 1.865 4.175 2.095 ;
        RECT 3.090 1.490 3.320 1.865 ;
        RECT 4.405 1.595 4.635 3.890 ;
        RECT 5.730 3.310 8.310 3.650 ;
        RECT 8.080 2.620 8.310 3.310 ;
        RECT 8.585 3.080 8.815 3.890 ;
        RECT 10.165 3.080 10.395 4.120 ;
        RECT 12.405 3.080 12.635 4.120 ;
        RECT 14.645 3.080 14.875 4.120 ;
        RECT 17.065 3.080 17.295 4.120 ;
        RECT 8.585 2.850 17.295 3.080 ;
        RECT 17.065 2.735 17.295 2.850 ;
        RECT 8.080 2.305 16.450 2.620 ;
        RECT 17.065 2.505 33.700 2.735 ;
        RECT 8.080 1.600 8.310 2.305 ;
        RECT 18.610 2.075 33.730 2.095 ;
        RECT 0.245 0.680 0.475 1.390 ;
        RECT 2.485 1.135 3.320 1.490 ;
        RECT 3.550 1.365 4.635 1.595 ;
        RECT 5.730 1.370 8.310 1.600 ;
        RECT 10.270 1.865 33.730 2.075 ;
        RECT 10.270 1.750 18.800 1.865 ;
        RECT 10.270 1.135 10.500 1.750 ;
        RECT 2.485 0.905 10.500 1.135 ;
        RECT 2.485 0.680 2.715 0.905 ;
        RECT 10.265 0.680 10.500 0.905 ;
        RECT 12.505 0.680 12.735 1.750 ;
        RECT 14.745 0.680 14.975 1.750 ;
        RECT 17.165 0.680 17.395 1.750 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_16
MACRO gf180mcu_fd_sc_mcu9t5v0__latq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.200 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.065 1.210 4.330 2.150 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.575 1.015 2.710 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.605 0.680 9.930 4.080 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 11.200 5.490 ;
        RECT 1.365 3.270 1.595 4.590 ;
        RECT 3.485 3.270 3.715 4.590 ;
        RECT 7.465 3.270 7.695 4.590 ;
        RECT 10.625 3.270 10.855 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 11.630 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 11.630 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.895 ;
        RECT 3.385 0.450 3.615 1.020 ;
        RECT 7.765 0.450 7.995 0.885 ;
        RECT 10.725 0.450 10.955 1.490 ;
        RECT 0.000 -0.450 11.200 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.270 0.575 4.080 ;
        RECT 0.245 1.345 0.475 3.270 ;
        RECT 2.665 2.610 2.895 4.080 ;
        RECT 5.245 3.410 5.475 4.080 ;
        RECT 5.245 3.180 6.215 3.410 ;
        RECT 5.525 2.610 5.755 2.950 ;
        RECT 2.665 2.380 5.755 2.610 ;
        RECT 2.085 1.355 2.315 1.915 ;
        RECT 1.085 1.345 2.315 1.355 ;
        RECT 0.245 1.125 2.315 1.345 ;
        RECT 0.245 1.115 1.155 1.125 ;
        RECT 0.245 0.680 0.475 1.115 ;
        RECT 2.665 0.680 2.895 2.380 ;
        RECT 4.665 1.575 4.895 2.380 ;
        RECT 5.985 1.345 6.215 3.180 ;
        RECT 8.485 2.375 8.735 4.080 ;
        RECT 7.085 2.365 8.735 2.375 ;
        RECT 7.085 2.145 9.115 2.365 ;
        RECT 7.085 1.575 7.315 2.145 ;
        RECT 8.205 1.345 8.435 1.915 ;
        RECT 5.985 1.225 8.435 1.345 ;
        RECT 5.345 1.115 8.435 1.225 ;
        RECT 5.345 0.885 6.190 1.115 ;
        RECT 8.665 0.975 9.115 2.145 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latq_1
MACRO gf180mcu_fd_sc_mcu9t5v0__latq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.320 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.065 1.210 4.330 2.150 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.575 1.015 2.710 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.675 1.590 11.050 4.235 ;
        RECT 10.230 1.210 11.050 1.590 ;
        RECT 10.725 0.680 11.050 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 12.320 5.490 ;
        RECT 1.365 3.425 1.595 4.590 ;
        RECT 3.485 3.425 3.715 4.590 ;
        RECT 7.465 3.425 7.695 4.590 ;
        RECT 9.655 3.425 9.885 4.590 ;
        RECT 11.695 3.425 11.925 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 12.750 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.750 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.895 ;
        RECT 3.385 0.450 3.615 1.020 ;
        RECT 7.765 0.450 7.995 0.885 ;
        RECT 9.605 0.450 9.835 1.490 ;
        RECT 11.845 0.450 12.075 1.490 ;
        RECT 0.000 -0.450 12.320 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.425 0.575 4.235 ;
        RECT 0.245 1.345 0.475 3.425 ;
        RECT 2.665 2.610 2.895 4.235 ;
        RECT 5.245 3.410 5.475 4.235 ;
        RECT 5.245 3.180 6.215 3.410 ;
        RECT 5.525 2.610 5.755 2.950 ;
        RECT 2.665 2.380 5.755 2.610 ;
        RECT 2.085 1.355 2.315 1.915 ;
        RECT 1.085 1.345 2.315 1.355 ;
        RECT 0.245 1.125 2.315 1.345 ;
        RECT 0.245 1.115 1.155 1.125 ;
        RECT 0.245 0.680 0.475 1.115 ;
        RECT 2.665 0.680 2.895 2.380 ;
        RECT 4.665 1.575 4.895 2.380 ;
        RECT 5.985 1.345 6.215 3.180 ;
        RECT 8.485 2.375 8.735 4.235 ;
        RECT 7.085 2.365 8.735 2.375 ;
        RECT 7.085 2.145 9.115 2.365 ;
        RECT 7.085 1.575 7.315 2.145 ;
        RECT 8.205 1.345 8.435 1.915 ;
        RECT 5.985 1.315 8.435 1.345 ;
        RECT 5.345 1.115 8.435 1.315 ;
        RECT 5.345 0.975 6.100 1.115 ;
        RECT 8.665 0.975 9.115 2.145 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latq_2
MACRO gf180mcu_fd_sc_mcu9t5v0__latq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.680 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.070 1.210 4.330 2.150 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 1.020 2.710 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.010 2.150 11.240 4.065 ;
        RECT 11.010 1.920 11.610 2.150 ;
        RECT 11.310 1.440 11.610 1.920 ;
        RECT 13.050 1.490 13.280 4.065 ;
        RECT 13.050 1.440 13.780 1.490 ;
        RECT 11.310 1.210 13.780 1.440 ;
        RECT 11.310 0.680 11.540 1.210 ;
        RECT 13.550 0.680 13.780 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 15.680 5.490 ;
        RECT 1.370 3.255 1.600 4.590 ;
        RECT 3.790 3.255 4.020 4.590 ;
        RECT 7.770 3.255 8.000 4.590 ;
        RECT 9.810 3.255 10.040 4.590 ;
        RECT 12.030 3.255 12.260 4.590 ;
        RECT 14.070 3.255 14.300 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 16.110 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 16.110 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.370 0.450 1.600 1.020 ;
        RECT 3.390 0.450 3.620 1.020 ;
        RECT 7.770 0.450 8.000 1.020 ;
        RECT 10.010 0.450 10.240 1.020 ;
        RECT 12.430 0.450 12.660 0.980 ;
        RECT 14.670 0.450 14.900 1.490 ;
        RECT 0.000 -0.450 15.680 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.250 3.255 0.580 4.065 ;
        RECT 0.250 1.540 0.480 3.255 ;
        RECT 2.570 2.720 2.800 4.065 ;
        RECT 5.550 3.180 5.780 4.065 ;
        RECT 5.550 2.950 6.520 3.180 ;
        RECT 2.570 2.380 6.060 2.720 ;
        RECT 1.990 1.540 2.220 2.150 ;
        RECT 0.250 1.310 2.220 1.540 ;
        RECT 0.250 0.680 0.480 1.310 ;
        RECT 2.570 0.680 2.900 2.380 ;
        RECT 4.670 1.810 4.900 2.380 ;
        RECT 6.290 1.020 6.520 2.950 ;
        RECT 8.790 2.610 9.120 4.065 ;
        RECT 7.330 2.380 9.120 2.610 ;
        RECT 7.330 1.810 7.560 2.380 ;
        RECT 8.210 1.480 8.440 2.150 ;
        RECT 5.350 0.910 6.520 1.020 ;
        RECT 7.310 1.250 8.440 1.480 ;
        RECT 7.310 0.910 7.540 1.250 ;
        RECT 5.350 0.680 7.540 0.910 ;
        RECT 8.890 0.680 9.120 2.380 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latq_4
MACRO gf180mcu_fd_sc_mcu9t5v0__latrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.880 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 1.770 3.295 2.710 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.084000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.965 2.440 5.500 2.670 ;
        RECT 0.705 1.540 0.970 2.295 ;
        RECT 3.675 1.725 4.135 2.295 ;
        RECT 4.965 1.725 5.195 2.440 ;
        RECT 3.675 1.540 5.195 1.725 ;
        RECT 0.705 1.495 5.195 1.540 ;
        RECT 0.705 1.310 3.905 1.495 ;
        RECT 0.705 1.210 0.970 1.310 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.340000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.455 2.710 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.910 0.845 12.355 4.360 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 12.880 5.490 ;
        RECT 1.265 3.550 1.495 4.590 ;
        RECT 3.025 3.860 3.255 4.590 ;
        RECT 6.630 3.550 6.860 4.590 ;
        RECT 9.215 3.550 9.445 4.590 ;
        RECT 11.055 3.875 11.285 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 13.310 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.310 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.080 ;
        RECT 7.145 0.450 7.375 1.135 ;
        RECT 9.165 0.450 9.395 1.135 ;
        RECT 11.005 0.450 11.235 1.605 ;
        RECT 0.000 -0.450 12.880 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.170 0.475 4.360 ;
        RECT 2.005 3.630 2.235 4.360 ;
        RECT 4.785 4.130 5.960 4.360 ;
        RECT 4.785 3.630 5.015 4.130 ;
        RECT 2.005 3.400 5.015 3.630 ;
        RECT 0.245 2.940 4.735 3.170 ;
        RECT 0.245 0.795 0.475 2.940 ;
        RECT 4.505 1.955 4.735 2.940 ;
        RECT 5.730 1.725 5.960 4.130 ;
        RECT 7.830 2.755 8.240 4.360 ;
        RECT 6.190 2.525 8.240 2.755 ;
        RECT 6.190 1.955 6.420 2.525 ;
        RECT 8.010 2.295 8.240 2.525 ;
        RECT 7.550 1.765 7.780 2.295 ;
        RECT 8.010 2.065 9.835 2.295 ;
        RECT 6.550 1.725 7.780 1.765 ;
        RECT 5.730 1.535 7.780 1.725 ;
        RECT 8.445 1.955 9.835 2.065 ;
        RECT 10.235 2.260 10.465 4.360 ;
        RECT 10.235 2.030 11.620 2.260 ;
        RECT 5.730 1.495 6.680 1.535 ;
        RECT 6.450 1.135 6.680 1.495 ;
        RECT 4.345 0.795 6.680 1.135 ;
        RECT 8.445 0.795 8.675 1.955 ;
        RECT 10.235 1.225 10.515 2.030 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrnq_1
MACRO gf180mcu_fd_sc_mcu9t5v0__latrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.000 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 1.770 3.260 2.710 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.084000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.770 2.765 5.380 2.995 ;
        RECT 4.770 2.150 5.000 2.765 ;
        RECT 0.895 1.835 1.600 2.065 ;
        RECT 1.370 1.540 1.600 1.835 ;
        RECT 4.070 1.780 5.000 2.150 ;
        RECT 4.070 1.540 4.330 1.780 ;
        RECT 1.370 1.310 4.330 1.540 ;
        RECT 4.070 1.210 4.330 1.310 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.340000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.065 2.090 2.710 ;
        RECT 1.830 1.770 2.475 2.065 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.355 0.845 12.730 4.360 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.000 5.490 ;
        RECT 1.390 3.550 1.620 4.590 ;
        RECT 3.130 3.860 3.360 4.590 ;
        RECT 6.650 3.690 6.880 4.590 ;
        RECT 9.420 3.550 9.650 4.590 ;
        RECT 11.335 3.880 11.565 4.590 ;
        RECT 13.375 3.880 13.605 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.430 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.430 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.435 0.450 1.775 1.080 ;
        RECT 7.350 0.450 7.580 1.135 ;
        RECT 9.370 0.450 9.600 1.135 ;
        RECT 11.285 0.450 11.515 1.605 ;
        RECT 13.525 0.450 13.755 1.605 ;
        RECT 0.000 -0.450 14.000 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.370 3.170 0.600 4.360 ;
        RECT 2.110 3.630 2.340 4.030 ;
        RECT 4.890 3.800 5.840 4.030 ;
        RECT 4.890 3.630 5.120 3.800 ;
        RECT 2.110 3.400 5.120 3.630 ;
        RECT 0.370 2.940 4.540 3.170 ;
        RECT 0.370 0.795 0.600 2.940 ;
        RECT 4.310 2.380 4.540 2.940 ;
        RECT 5.610 1.135 5.840 3.800 ;
        RECT 7.895 2.580 8.440 4.360 ;
        RECT 7.290 2.350 8.440 2.580 ;
        RECT 7.290 2.120 7.520 2.350 ;
        RECT 8.210 2.120 8.440 2.350 ;
        RECT 6.070 1.890 7.520 2.120 ;
        RECT 6.070 1.780 6.300 1.890 ;
        RECT 7.750 1.595 7.980 2.120 ;
        RECT 4.550 1.025 5.840 1.135 ;
        RECT 6.440 1.365 7.980 1.595 ;
        RECT 8.210 1.780 10.040 2.120 ;
        RECT 10.440 2.065 10.670 4.360 ;
        RECT 10.440 1.835 12.010 2.065 ;
        RECT 6.440 1.025 6.670 1.365 ;
        RECT 4.550 0.795 6.670 1.025 ;
        RECT 8.210 0.795 8.880 1.780 ;
        RECT 10.440 1.225 10.720 1.835 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrnq_2
MACRO gf180mcu_fd_sc_mcu9t5v0__latrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.500 1.770 3.770 2.720 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.084000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.740 1.540 0.970 2.720 ;
        RECT 4.120 1.585 4.350 2.720 ;
        RECT 5.640 2.150 5.870 2.720 ;
        RECT 5.190 1.920 5.870 2.150 ;
        RECT 5.190 1.585 5.450 1.920 ;
        RECT 4.120 1.540 5.450 1.585 ;
        RECT 0.740 1.355 5.450 1.540 ;
        RECT 0.740 1.310 4.260 1.355 ;
        RECT 5.190 1.210 5.450 1.355 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.340000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.390 1.770 2.650 2.720 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.035 3.645 14.265 4.360 ;
        RECT 16.075 3.645 16.305 4.360 ;
        RECT 14.035 3.415 16.305 3.645 ;
        RECT 14.035 2.055 14.410 3.415 ;
        RECT 14.035 1.825 16.555 2.055 ;
        RECT 14.035 0.785 14.410 1.825 ;
        RECT 16.325 0.785 16.555 1.825 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.920 5.490 ;
        RECT 1.320 3.550 1.550 4.590 ;
        RECT 3.240 3.870 3.470 4.590 ;
        RECT 7.610 3.700 7.840 4.590 ;
        RECT 9.880 3.550 10.110 4.590 ;
        RECT 12.070 3.550 12.300 4.590 ;
        RECT 13.015 3.875 13.245 4.590 ;
        RECT 15.055 3.875 15.285 4.590 ;
        RECT 17.095 3.875 17.325 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 18.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.345 0.450 1.685 1.070 ;
        RECT 7.740 0.450 7.970 1.125 ;
        RECT 9.980 0.450 10.210 1.125 ;
        RECT 12.220 0.450 12.450 1.125 ;
        RECT 12.965 0.450 13.195 1.595 ;
        RECT 15.205 0.450 15.435 1.595 ;
        RECT 17.445 0.450 17.675 1.595 ;
        RECT 0.000 -0.450 17.920 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.280 3.180 0.530 4.360 ;
        RECT 2.220 3.640 2.450 4.040 ;
        RECT 5.320 3.810 6.330 4.040 ;
        RECT 5.320 3.640 5.550 3.810 ;
        RECT 2.220 3.410 5.550 3.640 ;
        RECT 0.280 2.950 5.270 3.180 ;
        RECT 0.280 0.785 0.510 2.950 ;
        RECT 5.040 2.380 5.270 2.950 ;
        RECT 6.100 2.150 6.330 3.810 ;
        RECT 8.810 3.180 9.040 4.360 ;
        RECT 11.050 3.550 11.325 4.360 ;
        RECT 7.170 2.950 10.840 3.180 ;
        RECT 7.170 2.380 7.400 2.950 ;
        RECT 8.230 2.150 8.460 2.720 ;
        RECT 6.100 1.920 8.460 2.150 ;
        RECT 4.580 0.980 4.810 1.125 ;
        RECT 6.100 0.980 6.330 1.920 ;
        RECT 4.580 0.750 6.330 0.980 ;
        RECT 8.860 0.785 9.090 2.950 ;
        RECT 10.610 2.380 10.840 2.950 ;
        RECT 11.095 2.665 11.325 3.550 ;
        RECT 11.095 2.435 13.740 2.665 ;
        RECT 11.095 0.785 11.330 2.435 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrnq_4
MACRO gf180mcu_fd_sc_mcu9t5v0__latrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.440 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 1.770 3.335 2.710 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.084000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 2.275 1.600 2.505 ;
        RECT 1.370 1.540 1.600 2.275 ;
        RECT 3.945 2.150 4.175 2.560 ;
        RECT 5.265 2.150 5.495 2.560 ;
        RECT 3.945 1.770 5.495 2.150 ;
        RECT 3.945 1.540 4.175 1.770 ;
        RECT 1.370 1.310 4.175 1.540 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.340000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.495 2.710 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.550 1.770 8.875 2.710 ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.425 0.845 12.735 4.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 13.440 5.490 ;
        RECT 1.265 3.400 1.495 4.590 ;
        RECT 3.065 3.890 3.295 4.590 ;
        RECT 6.645 3.890 6.875 4.590 ;
        RECT 8.925 3.400 9.155 4.590 ;
        RECT 11.225 3.430 11.455 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 13.870 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.870 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.080 ;
        RECT 7.130 0.450 7.470 1.075 ;
        RECT 11.385 0.450 11.615 1.165 ;
        RECT 0.000 -0.450 13.440 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.170 0.475 4.210 ;
        RECT 2.045 3.630 2.275 4.210 ;
        RECT 4.825 3.630 5.055 4.210 ;
        RECT 2.045 3.400 7.315 3.630 ;
        RECT 0.245 2.940 4.775 3.170 ;
        RECT 7.085 3.020 7.315 3.400 ;
        RECT 0.245 0.790 0.475 2.940 ;
        RECT 4.545 2.380 4.775 2.940 ;
        RECT 5.725 2.790 7.315 3.020 ;
        RECT 7.905 3.170 8.135 4.210 ;
        RECT 10.205 3.200 10.435 4.210 ;
        RECT 7.905 2.940 9.555 3.170 ;
        RECT 10.205 2.970 11.915 3.200 ;
        RECT 5.725 1.130 5.955 2.790 ;
        RECT 9.325 2.560 9.555 2.940 ;
        RECT 6.185 1.540 6.415 2.560 ;
        RECT 9.325 2.220 10.715 2.560 ;
        RECT 9.325 1.540 9.555 2.220 ;
        RECT 11.685 1.655 11.915 2.970 ;
        RECT 6.185 1.310 9.555 1.540 ;
        RECT 10.045 1.425 11.915 1.655 ;
        RECT 10.045 1.315 10.275 1.425 ;
        RECT 4.385 0.790 5.955 1.130 ;
        RECT 9.325 0.790 9.555 1.310 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrsnq_1
MACRO gf180mcu_fd_sc_mcu9t5v0__latrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.020000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 2.505 3.210 3.270 ;
        RECT 2.950 2.275 3.810 2.505 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.322000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.925 1.990 1.155 2.560 ;
        RECT 4.070 1.990 4.755 2.710 ;
        RECT 5.885 1.990 6.115 2.560 ;
        RECT 0.925 1.760 6.115 1.990 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.440000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.275 2.650 2.710 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.302000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.110 1.770 9.535 2.710 ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.945 2.150 13.175 4.310 ;
        RECT 12.470 1.210 13.175 2.150 ;
        RECT 12.945 0.790 13.175 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.560 5.490 ;
        RECT 1.365 3.880 1.595 4.590 ;
        RECT 3.425 4.420 3.655 4.590 ;
        RECT 7.565 3.500 7.795 4.590 ;
        RECT 9.985 3.880 10.215 4.590 ;
        RECT 11.825 3.880 12.055 4.590 ;
        RECT 14.065 3.880 14.295 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.585 0.450 1.815 1.130 ;
        RECT 7.605 0.450 7.835 1.130 ;
        RECT 11.825 0.450 12.055 1.530 ;
        RECT 14.065 0.450 14.295 1.600 ;
        RECT 0.000 -0.450 14.560 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.650 0.475 4.310 ;
        RECT 2.085 4.190 2.315 4.220 ;
        RECT 5.605 4.190 5.835 4.310 ;
        RECT 2.085 3.960 5.835 4.190 ;
        RECT 2.085 3.880 2.315 3.960 ;
        RECT 2.490 3.650 5.355 3.730 ;
        RECT 0.245 3.500 5.355 3.650 ;
        RECT 0.245 3.420 2.665 3.500 ;
        RECT 0.245 0.790 0.695 3.420 ;
        RECT 5.125 2.220 5.355 3.500 ;
        RECT 5.605 3.020 5.835 3.960 ;
        RECT 8.865 3.650 9.095 4.310 ;
        RECT 10.705 3.650 10.935 4.310 ;
        RECT 8.865 3.420 9.995 3.650 ;
        RECT 10.705 3.420 12.240 3.650 ;
        RECT 5.605 2.790 8.235 3.020 ;
        RECT 6.345 1.130 6.575 2.790 ;
        RECT 7.135 1.990 7.365 2.560 ;
        RECT 8.005 2.220 8.235 2.790 ;
        RECT 9.765 2.560 9.995 3.420 ;
        RECT 9.765 2.220 11.375 2.560 ;
        RECT 7.135 1.760 8.210 1.990 ;
        RECT 7.980 1.540 8.210 1.760 ;
        RECT 9.765 1.540 9.995 2.220 ;
        RECT 12.010 1.990 12.240 3.420 ;
        RECT 7.980 1.310 9.995 1.540 ;
        RECT 4.805 0.790 6.575 1.130 ;
        RECT 9.745 0.790 9.995 1.310 ;
        RECT 10.705 1.760 12.240 1.990 ;
        RECT 10.705 0.790 10.935 1.760 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrsnq_2
MACRO gf180mcu_fd_sc_mcu9t5v0__latrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.360 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 2.195 3.210 2.710 ;
        RECT 2.950 1.770 3.500 2.195 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.084000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.525 2.875 5.370 3.105 ;
        RECT 1.830 2.195 2.090 2.710 ;
        RECT 0.970 1.965 2.090 2.195 ;
        RECT 4.525 2.120 4.755 2.875 ;
        RECT 1.830 1.540 2.090 1.965 ;
        RECT 4.055 1.890 4.755 2.120 ;
        RECT 4.055 1.540 4.285 1.890 ;
        RECT 1.830 1.310 4.285 1.540 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.340000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.375 1.770 2.650 2.710 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.550 1.770 8.985 2.710 ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.265 3.650 13.495 4.290 ;
        RECT 15.305 3.650 15.535 4.290 ;
        RECT 13.265 3.420 15.535 3.650 ;
        RECT 13.515 2.150 13.745 3.420 ;
        RECT 13.515 1.920 15.530 2.150 ;
        RECT 13.515 0.845 13.745 1.920 ;
        RECT 15.270 1.655 15.530 1.920 ;
        RECT 15.270 1.210 15.985 1.655 ;
        RECT 15.755 0.845 15.985 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.360 5.490 ;
        RECT 1.305 3.480 1.535 4.590 ;
        RECT 3.045 4.120 3.275 4.590 ;
        RECT 6.565 3.480 6.795 4.590 ;
        RECT 8.785 3.650 9.015 4.590 ;
        RECT 10.205 3.880 10.435 4.590 ;
        RECT 12.245 3.880 12.475 4.590 ;
        RECT 14.285 3.880 14.515 4.590 ;
        RECT 16.325 3.880 16.555 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 17.790 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 17.790 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.460 0.450 1.800 1.080 ;
        RECT 7.240 0.450 7.580 1.080 ;
        RECT 10.155 0.450 10.385 1.165 ;
        RECT 12.395 0.450 12.625 1.165 ;
        RECT 14.635 0.450 14.865 1.165 ;
        RECT 16.875 0.450 17.105 1.165 ;
        RECT 0.000 -0.450 17.360 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.285 3.170 0.515 4.290 ;
        RECT 2.025 3.710 2.255 4.290 ;
        RECT 4.805 3.710 5.035 4.290 ;
        RECT 2.025 3.565 5.035 3.710 ;
        RECT 2.025 3.480 5.830 3.565 ;
        RECT 4.820 3.335 5.830 3.480 ;
        RECT 0.285 2.940 4.295 3.170 ;
        RECT 0.285 0.795 0.625 2.940 ;
        RECT 4.065 2.380 4.295 2.940 ;
        RECT 5.600 2.720 5.830 3.335 ;
        RECT 7.765 3.420 7.995 4.290 ;
        RECT 7.765 3.190 9.665 3.420 ;
        RECT 5.600 2.655 7.535 2.720 ;
        RECT 5.535 2.490 7.535 2.655 ;
        RECT 5.535 1.135 5.765 2.490 ;
        RECT 6.135 1.540 6.365 2.260 ;
        RECT 7.305 1.935 7.535 2.490 ;
        RECT 9.435 2.250 9.665 3.190 ;
        RECT 11.225 2.760 11.455 4.290 ;
        RECT 11.225 2.530 12.915 2.760 ;
        RECT 9.435 1.910 11.065 2.250 ;
        RECT 9.435 1.540 9.665 1.910 ;
        RECT 12.685 1.655 12.915 2.530 ;
        RECT 6.135 1.310 9.665 1.540 ;
        RECT 4.495 0.795 5.765 1.135 ;
        RECT 9.435 0.795 9.665 1.310 ;
        RECT 11.275 1.425 12.915 1.655 ;
        RECT 11.275 0.845 11.505 1.425 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrsnq_4
MACRO gf180mcu_fd_sc_mcu9t5v0__latsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.760 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.210 2.270 2.160 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.084000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.390 3.295 2.620 ;
        RECT 0.710 1.770 1.015 2.390 ;
        RECT 3.065 2.090 3.295 2.390 ;
        RECT 3.690 2.090 4.030 3.200 ;
        RECT 3.065 1.830 4.030 2.090 ;
    END
  END E
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.870 1.210 7.210 2.160 ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.720 0.845 11.050 4.230 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 11.760 5.490 ;
        RECT 1.365 3.420 1.595 4.590 ;
        RECT 5.225 3.420 5.455 4.590 ;
        RECT 7.685 3.420 7.915 4.590 ;
        RECT 9.570 3.420 9.800 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 12.190 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.190 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.185 ;
        RECT 5.465 0.450 5.695 1.185 ;
        RECT 9.700 0.450 9.930 1.220 ;
        RECT 0.000 -0.450 11.760 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.190 0.575 4.230 ;
        RECT 3.305 4.000 4.490 4.230 ;
        RECT 3.305 3.420 3.535 4.000 ;
        RECT 0.245 2.850 2.955 3.190 ;
        RECT 0.245 0.845 0.475 2.850 ;
        RECT 4.260 1.185 4.490 4.000 ;
        RECT 6.665 2.675 6.895 4.230 ;
        RECT 8.500 3.205 8.730 4.230 ;
        RECT 8.500 2.975 9.485 3.205 ;
        RECT 5.625 2.620 6.895 2.675 ;
        RECT 5.625 2.445 7.835 2.620 ;
        RECT 5.625 2.215 5.855 2.445 ;
        RECT 6.745 2.390 7.835 2.445 ;
        RECT 7.605 2.215 7.835 2.390 ;
        RECT 4.785 1.875 5.855 2.215 ;
        RECT 6.085 1.645 6.315 2.215 ;
        RECT 3.505 1.075 4.490 1.185 ;
        RECT 5.005 1.415 6.315 1.645 ;
        RECT 7.605 1.875 9.025 2.215 ;
        RECT 9.255 1.935 9.485 2.975 ;
        RECT 10.140 1.935 10.370 2.215 ;
        RECT 5.005 1.075 5.235 1.415 ;
        RECT 3.505 0.845 5.235 1.075 ;
        RECT 7.605 0.845 7.835 1.875 ;
        RECT 9.255 1.790 10.370 1.935 ;
        RECT 9.240 1.705 10.370 1.790 ;
        RECT 9.240 1.225 9.470 1.705 ;
        RECT 8.355 0.885 9.470 1.225 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latsnq_1
MACRO gf180mcu_fd_sc_mcu9t5v0__latsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.320 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.210 2.090 2.335 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.084000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.235 3.090 4.080 3.320 ;
        RECT 3.235 2.795 3.465 3.090 ;
        RECT 0.925 2.565 3.465 2.795 ;
        RECT 0.925 1.995 1.155 2.565 ;
        RECT 2.950 2.050 3.465 2.565 ;
        RECT 2.950 1.770 3.210 2.050 ;
    END
  END E
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.870 1.770 7.155 2.710 ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.575 2.150 10.805 4.200 ;
        RECT 10.575 0.680 11.050 2.150 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 12.320 5.490 ;
        RECT 1.415 3.665 1.645 4.590 ;
        RECT 5.115 3.550 5.345 4.590 ;
        RECT 7.335 3.550 7.565 4.590 ;
        RECT 9.555 3.860 9.785 4.590 ;
        RECT 11.595 3.550 11.825 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 12.750 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.750 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.020 ;
        RECT 5.465 0.450 5.695 1.020 ;
        RECT 9.605 0.450 9.835 1.305 ;
        RECT 11.845 0.450 12.075 1.490 ;
        RECT 0.000 -0.450 12.320 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.365 0.625 4.360 ;
        RECT 3.355 4.130 4.540 4.360 ;
        RECT 3.355 3.550 3.585 4.130 ;
        RECT 0.245 3.025 3.005 3.365 ;
        RECT 0.245 0.680 0.475 3.025 ;
        RECT 4.310 1.765 4.540 4.130 ;
        RECT 6.315 3.170 6.545 4.200 ;
        RECT 8.535 3.630 8.765 4.210 ;
        RECT 8.535 3.400 10.225 3.630 ;
        RECT 5.025 2.940 9.205 3.170 ;
        RECT 5.025 1.995 5.255 2.940 ;
        RECT 5.735 1.765 5.965 2.335 ;
        RECT 8.975 2.225 9.205 2.940 ;
        RECT 3.505 1.535 5.965 1.765 ;
        RECT 7.605 1.995 9.205 2.225 ;
        RECT 3.505 0.680 3.735 1.535 ;
        RECT 7.605 0.680 7.835 1.995 ;
        RECT 9.995 1.765 10.225 3.400 ;
        RECT 8.485 1.535 10.225 1.765 ;
        RECT 8.485 0.680 8.715 1.535 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latsnq_2
MACRO gf180mcu_fd_sc_mcu9t5v0__latsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.680 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.245 1.210 2.650 2.150 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 2.084000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 2.945 4.195 3.270 ;
        RECT 3.510 2.610 3.770 2.945 ;
        RECT 1.785 2.380 3.770 2.610 ;
        RECT 1.785 2.150 2.015 2.380 ;
        RECT 0.945 1.920 2.015 2.150 ;
        RECT 2.880 2.330 3.770 2.380 ;
        RECT 2.880 1.920 3.220 2.330 ;
    END
  END E
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.870 1.770 7.230 2.710 ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.510 3.320 11.740 4.250 ;
        RECT 13.550 3.320 13.780 4.250 ;
        RECT 11.510 3.090 13.780 3.320 ;
        RECT 11.760 1.440 11.990 3.090 ;
        RECT 13.590 1.650 13.850 2.150 ;
        RECT 13.590 1.440 14.230 1.650 ;
        RECT 11.760 1.210 14.230 1.440 ;
        RECT 11.760 0.840 11.990 1.210 ;
        RECT 14.000 0.840 14.230 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 15.680 5.490 ;
        RECT 1.610 3.705 1.840 4.590 ;
        RECT 5.390 3.550 5.620 4.590 ;
        RECT 7.610 3.875 7.840 4.590 ;
        RECT 8.450 3.875 8.680 4.590 ;
        RECT 10.490 3.875 10.720 4.590 ;
        RECT 12.530 3.550 12.760 4.590 ;
        RECT 14.570 3.875 14.800 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 16.110 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 16.110 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.440 0.450 1.670 1.305 ;
        RECT 5.540 0.450 5.770 1.310 ;
        RECT 8.400 0.450 8.630 1.160 ;
        RECT 10.640 0.450 10.870 1.160 ;
        RECT 12.880 0.450 13.110 0.690 ;
        RECT 15.120 0.450 15.350 1.160 ;
        RECT 0.000 -0.450 15.680 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.590 3.180 0.820 4.360 ;
        RECT 3.630 4.130 4.655 4.360 ;
        RECT 3.630 3.550 3.860 4.130 ;
        RECT 0.590 2.890 3.280 3.180 ;
        RECT 0.320 2.840 3.280 2.890 ;
        RECT 0.320 2.660 0.815 2.840 ;
        RECT 0.320 0.880 0.550 2.660 ;
        RECT 4.425 1.770 4.655 4.130 ;
        RECT 6.590 3.170 6.820 4.250 ;
        RECT 6.590 3.135 9.070 3.170 ;
        RECT 5.100 2.940 9.070 3.135 ;
        RECT 5.100 2.905 6.715 2.940 ;
        RECT 5.100 2.000 5.330 2.905 ;
        RECT 6.000 1.770 6.230 2.310 ;
        RECT 3.580 1.540 6.230 1.770 ;
        RECT 8.840 1.650 9.070 2.940 ;
        RECT 3.580 0.970 3.810 1.540 ;
        RECT 7.680 1.420 9.070 1.650 ;
        RECT 9.470 2.280 9.700 4.250 ;
        RECT 9.470 1.940 11.300 2.280 ;
        RECT 7.680 0.840 7.910 1.420 ;
        RECT 9.470 0.840 9.750 1.940 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latsnq_4
MACRO gf180mcu_fd_sc_mcu9t5v0__mux2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.853500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.630 1.770 5.450 2.150 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.853500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.390 1.770 2.650 2.710 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 2.705 6.035 3.270 ;
        RECT 3.225 2.475 6.035 2.705 ;
        RECT 3.225 1.380 3.455 2.475 ;
        RECT 5.750 1.770 6.035 2.475 ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 0.720 0.575 4.235 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.280 5.490 ;
        RECT 1.365 2.970 1.595 4.590 ;
        RECT 5.310 3.480 5.650 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.060 ;
        RECT 5.465 0.450 5.695 0.990 ;
        RECT 0.000 -0.450 7.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.930 3.545 3.835 3.775 ;
        RECT 1.930 2.055 2.160 3.545 ;
        RECT 3.605 2.965 3.835 3.545 ;
        RECT 0.870 1.825 2.160 2.055 ;
        RECT 1.930 1.005 2.160 1.825 ;
        RECT 3.945 1.540 4.175 2.110 ;
        RECT 6.385 1.540 6.815 3.775 ;
        RECT 3.945 1.310 6.815 1.540 ;
        RECT 1.930 0.775 3.790 1.005 ;
        RECT 6.585 0.720 6.815 1.310 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux2_1
MACRO gf180mcu_fd_sc_mcu9t5v0__mux2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.400 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 1.770 6.570 2.150 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 1.770 3.255 2.710 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.005 2.470 7.315 2.710 ;
        RECT 4.005 1.775 4.235 2.470 ;
        RECT 6.870 1.770 7.315 2.470 ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.729500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 0.680 1.595 4.360 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 8.400 5.490 ;
        RECT 0.295 3.550 0.525 4.590 ;
        RECT 2.385 3.550 2.615 4.590 ;
        RECT 6.645 3.550 6.875 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 8.830 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.830 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.020 ;
        RECT 6.645 0.450 6.875 1.020 ;
        RECT 0.000 -0.450 8.400 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 4.885 3.170 5.115 4.360 ;
        RECT 1.945 2.940 5.115 3.170 ;
        RECT 1.945 1.540 2.175 2.940 ;
        RECT 4.830 1.830 5.520 2.060 ;
        RECT 5.290 1.540 5.520 1.830 ;
        RECT 7.665 1.540 7.995 4.360 ;
        RECT 1.945 1.310 4.675 1.540 ;
        RECT 5.290 1.310 7.995 1.540 ;
        RECT 4.445 0.680 4.675 1.310 ;
        RECT 7.765 0.680 7.995 1.310 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux2_2
MACRO gf180mcu_fd_sc_mcu9t5v0__mux2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.640 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.990 1.830 8.645 2.150 ;
        RECT 7.990 1.210 8.250 1.830 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.130 1.770 6.010 2.150 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.300 2.470 9.430 2.700 ;
        RECT 6.300 1.775 6.530 2.470 ;
        RECT 9.050 2.060 9.430 2.470 ;
        RECT 9.050 1.830 9.665 2.060 ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.550500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.420 2.710 1.650 4.360 ;
        RECT 3.610 2.710 3.890 4.360 ;
        RECT 1.420 2.330 3.890 2.710 ;
        RECT 1.420 0.680 1.650 2.330 ;
        RECT 3.660 0.680 3.890 2.330 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 10.640 5.490 ;
        RECT 0.350 3.550 0.580 4.590 ;
        RECT 2.490 3.550 2.720 4.590 ;
        RECT 4.680 3.550 4.910 4.590 ;
        RECT 8.940 3.550 9.170 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 11.070 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 11.070 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 0.450 0.530 1.490 ;
        RECT 2.540 0.450 2.770 1.490 ;
        RECT 4.780 0.450 5.010 1.020 ;
        RECT 8.940 0.450 9.170 1.020 ;
        RECT 0.000 -0.450 10.640 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 7.180 3.160 7.410 4.360 ;
        RECT 4.670 2.930 7.410 3.160 ;
        RECT 4.670 2.115 4.900 2.930 ;
        RECT 4.240 1.775 4.900 2.115 ;
        RECT 7.125 1.830 7.760 2.060 ;
        RECT 4.670 1.540 4.900 1.775 ;
        RECT 4.670 1.310 6.970 1.540 ;
        RECT 6.740 0.680 6.970 1.310 ;
        RECT 7.530 0.980 7.760 1.830 ;
        RECT 9.960 1.480 10.290 4.360 ;
        RECT 8.480 1.250 10.290 1.480 ;
        RECT 8.480 0.980 8.710 1.250 ;
        RECT 7.530 0.750 8.710 0.980 ;
        RECT 10.060 0.680 10.290 1.250 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux2_4
MACRO gf180mcu_fd_sc_mcu9t5v0__mux4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.360 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.853500 ;
    PORT
      LAYER Metal1 ;
        RECT 14.710 1.210 14.970 2.555 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.853500 ;
    PORT
      LAYER Metal1 ;
        RECT 11.350 1.770 11.610 2.710 ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.853500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 0.970 2.710 ;
    END
  END I2
  PIN I3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.853500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.070 1.770 4.375 2.710 ;
    END
  END I3
  PIN S0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.390 1.900 2.650 2.995 ;
        RECT 2.390 1.670 3.210 1.900 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.405 2.155 8.810 3.195 ;
        RECT 7.675 1.770 8.810 2.155 ;
    END
  END S1
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.003200 ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 2.330 6.255 3.175 ;
        RECT 6.025 1.590 6.255 2.330 ;
        RECT 5.750 1.210 6.255 1.590 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.360 5.490 ;
        RECT 0.295 3.440 0.525 4.590 ;
        RECT 4.725 3.865 4.955 4.590 ;
        RECT 10.935 3.440 11.165 4.590 ;
        RECT 15.015 3.440 15.245 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.280 17.790 5.470 ;
        RECT -0.430 2.265 0.430 2.280 ;
        RECT 16.930 2.265 17.790 2.280 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 4.745 2.265 6.455 2.280 ;
        RECT -0.430 -0.430 17.790 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.430 ;
        RECT 4.725 0.450 4.955 1.430 ;
        RECT 10.835 0.450 11.065 1.430 ;
        RECT 15.315 0.450 15.545 1.430 ;
        RECT 0.000 -0.450 17.360 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 1.090 1.595 4.170 ;
        RECT 2.665 3.940 4.495 4.170 ;
        RECT 2.665 3.455 2.895 3.940 ;
        RECT 1.930 3.225 2.895 3.455 ;
        RECT 3.605 3.355 3.915 3.695 ;
        RECT 4.265 3.635 4.495 3.940 ;
        RECT 6.805 3.635 7.035 4.170 ;
        RECT 4.265 3.405 7.035 3.635 ;
        RECT 6.755 3.360 7.035 3.405 ;
        RECT 1.930 1.375 2.160 3.225 ;
        RECT 1.930 1.145 2.770 1.375 ;
        RECT 3.605 1.090 3.835 3.355 ;
        RECT 5.290 1.790 5.575 2.130 ;
        RECT 5.290 0.925 5.520 1.790 ;
        RECT 6.755 1.155 6.985 3.360 ;
        RECT 7.825 2.615 8.055 4.170 ;
        RECT 8.845 4.005 10.705 4.235 ;
        RECT 8.845 3.425 9.270 4.005 ;
        RECT 7.215 2.385 8.055 2.615 ;
        RECT 7.215 0.925 7.445 2.385 ;
        RECT 9.040 1.430 9.270 3.425 ;
        RECT 9.915 2.315 10.145 3.695 ;
        RECT 10.475 3.210 10.705 4.005 ;
        RECT 11.395 3.940 13.305 4.170 ;
        RECT 11.395 3.210 11.625 3.940 ;
        RECT 10.475 2.980 11.625 3.210 ;
        RECT 7.875 0.925 8.105 1.345 ;
        RECT 8.995 1.090 9.270 1.430 ;
        RECT 9.500 1.090 10.145 2.315 ;
        RECT 11.955 1.090 12.185 3.695 ;
        RECT 12.975 1.090 13.305 3.940 ;
        RECT 13.995 3.475 14.225 4.250 ;
        RECT 13.675 3.245 14.225 3.475 ;
        RECT 13.675 1.375 13.905 3.245 ;
        RECT 16.035 3.015 16.265 4.170 ;
        RECT 14.135 2.785 16.665 3.015 ;
        RECT 14.135 2.215 14.365 2.785 ;
        RECT 13.675 1.145 14.480 1.375 ;
        RECT 16.435 1.090 16.665 2.785 ;
        RECT 5.290 0.695 8.105 0.925 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux4_1
MACRO gf180mcu_fd_sc_mcu9t5v0__mux4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.120000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.950 1.210 17.210 2.030 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.120000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.590 1.770 13.850 2.390 ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.120000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.050 1.015 3.270 ;
    END
  END I2
  PIN I3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.120000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.625 2.050 4.890 2.710 ;
    END
  END I3
  PIN S0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.360000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.285 2.000 2.515 2.390 ;
        RECT 3.510 2.000 3.815 2.260 ;
        RECT 2.285 1.770 3.815 2.000 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.240000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.600 2.150 10.830 2.830 ;
        RECT 9.560 1.770 10.830 2.150 ;
        RECT 9.560 1.690 9.790 1.770 ;
    END
  END S1
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.081600 ;
    PORT
      LAYER Metal1 ;
        RECT 6.310 1.200 6.755 3.380 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 19.040 5.490 ;
        RECT 0.250 3.080 0.480 4.590 ;
        RECT 5.285 4.070 5.515 4.590 ;
        RECT 7.545 3.080 7.775 4.590 ;
        RECT 13.000 3.080 13.230 4.590 ;
        RECT 17.340 3.080 17.570 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 19.470 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 19.470 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.540 ;
        RECT 5.405 0.450 5.635 1.540 ;
        RECT 7.645 0.450 7.875 1.540 ;
        RECT 12.960 0.450 13.190 1.540 ;
        RECT 17.440 0.450 17.670 1.540 ;
        RECT 0.000 -0.450 19.040 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 11.120 4.120 12.770 4.350 ;
        RECT 1.365 1.200 1.595 3.890 ;
        RECT 1.825 3.840 2.955 3.890 ;
        RECT 1.825 3.610 7.315 3.840 ;
        RECT 1.825 1.485 2.055 3.610 ;
        RECT 2.725 3.080 2.955 3.610 ;
        RECT 4.045 1.845 4.275 3.380 ;
        RECT 7.085 2.850 7.315 3.610 ;
        RECT 8.640 3.080 9.005 3.890 ;
        RECT 9.235 3.660 10.180 3.890 ;
        RECT 8.640 2.850 8.870 3.080 ;
        RECT 7.085 2.620 8.870 2.850 ;
        RECT 7.105 2.000 7.335 2.390 ;
        RECT 4.045 1.615 4.515 1.845 ;
        RECT 7.105 1.770 8.410 2.000 ;
        RECT 1.825 1.255 3.450 1.485 ;
        RECT 4.285 1.200 4.515 1.615 ;
        RECT 8.180 0.980 8.410 1.770 ;
        RECT 8.640 1.210 8.870 2.620 ;
        RECT 9.235 2.570 9.465 3.660 ;
        RECT 9.950 3.080 10.180 3.660 ;
        RECT 9.100 2.360 9.465 2.570 ;
        RECT 9.100 0.980 9.330 2.360 ;
        RECT 10.000 0.980 10.230 1.540 ;
        RECT 11.120 1.200 11.410 4.120 ;
        RECT 11.680 1.200 12.210 3.890 ;
        RECT 12.540 2.850 12.770 4.120 ;
        RECT 13.460 4.120 15.430 4.350 ;
        RECT 13.460 2.850 13.690 4.120 ;
        RECT 12.540 2.620 13.690 2.850 ;
        RECT 14.080 1.200 14.310 3.890 ;
        RECT 15.170 1.200 15.430 4.120 ;
        RECT 16.190 2.895 16.420 3.890 ;
        RECT 15.700 2.665 16.420 2.895 ;
        RECT 15.700 1.485 15.930 2.665 ;
        RECT 18.460 2.490 18.790 3.890 ;
        RECT 16.570 2.435 18.790 2.490 ;
        RECT 16.160 2.260 18.790 2.435 ;
        RECT 16.160 2.050 16.720 2.260 ;
        RECT 15.700 1.255 16.605 1.485 ;
        RECT 18.560 1.200 18.790 2.260 ;
        RECT 8.180 0.750 10.230 0.980 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux4_2
MACRO gf180mcu_fd_sc_mcu9t5v0__mux4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.120000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.190 1.210 19.450 2.030 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.120000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.830 2.150 16.090 2.710 ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.120000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.700 2.330 1.080 2.710 ;
    END
  END I2
  PIN I3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.120000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.630 2.150 4.890 2.710 ;
    END
  END I3
  PIN S0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.360000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.350 2.220 2.580 2.710 ;
        RECT 2.350 1.770 3.885 2.220 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.240000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.905 2.175 13.135 2.830 ;
        RECT 11.790 1.945 13.135 2.175 ;
        RECT 12.470 1.210 12.730 1.945 ;
    END
  END S1
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.163200 ;
    PORT
      LAYER Metal1 ;
        RECT 6.590 2.030 6.825 3.380 ;
        RECT 9.075 2.030 9.370 3.380 ;
        RECT 6.590 1.800 9.370 2.030 ;
        RECT 6.590 1.230 6.820 1.800 ;
        RECT 8.830 1.210 9.370 1.800 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 21.280 5.490 ;
        RECT 0.410 3.040 0.640 4.590 ;
        RECT 5.355 4.070 5.585 4.590 ;
        RECT 7.835 4.070 8.065 4.590 ;
        RECT 10.095 3.440 10.325 4.590 ;
        RECT 15.245 3.400 15.475 4.590 ;
        RECT 19.585 3.040 19.815 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 21.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.310 0.450 0.540 1.570 ;
        RECT 5.470 0.450 5.700 1.570 ;
        RECT 7.710 0.450 7.940 1.570 ;
        RECT 9.950 0.450 10.180 1.570 ;
        RECT 15.205 0.450 15.435 1.570 ;
        RECT 19.685 0.450 19.915 1.570 ;
        RECT 0.000 -0.450 21.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 13.465 4.080 15.015 4.310 ;
        RECT 1.430 1.230 1.660 3.850 ;
        RECT 1.890 3.840 3.020 3.850 ;
        RECT 1.890 3.610 9.865 3.840 ;
        RECT 1.890 1.515 2.120 3.610 ;
        RECT 2.790 3.040 3.020 3.610 ;
        RECT 4.115 1.925 4.345 3.380 ;
        RECT 9.635 3.210 9.865 3.610 ;
        RECT 11.425 3.270 11.655 3.850 ;
        RECT 10.945 3.210 11.655 3.270 ;
        RECT 9.635 3.040 11.655 3.210 ;
        RECT 9.635 2.980 11.100 3.040 ;
        RECT 9.655 2.030 9.885 2.710 ;
        RECT 4.115 1.695 4.580 1.925 ;
        RECT 9.655 1.800 10.640 2.030 ;
        RECT 1.890 1.285 3.515 1.515 ;
        RECT 4.350 1.230 4.580 1.695 ;
        RECT 10.410 1.000 10.640 1.800 ;
        RECT 10.870 1.230 11.100 2.980 ;
        RECT 12.445 2.635 12.675 3.850 ;
        RECT 11.330 2.405 12.675 2.635 ;
        RECT 11.330 1.000 11.560 2.405 ;
        RECT 13.465 1.570 13.695 4.080 ;
        RECT 12.005 1.000 12.235 1.570 ;
        RECT 13.125 1.230 13.695 1.570 ;
        RECT 13.925 1.230 14.455 3.850 ;
        RECT 14.785 3.170 15.015 4.080 ;
        RECT 15.705 4.080 17.675 4.310 ;
        RECT 15.705 3.170 15.935 4.080 ;
        RECT 14.785 2.940 15.935 3.170 ;
        RECT 16.325 1.230 16.555 3.850 ;
        RECT 17.445 1.230 17.675 4.080 ;
        RECT 18.565 2.950 18.795 3.850 ;
        RECT 17.945 2.720 18.795 2.950 ;
        RECT 17.945 1.515 18.175 2.720 ;
        RECT 20.705 2.490 21.035 3.850 ;
        RECT 18.405 2.260 21.035 2.490 ;
        RECT 18.405 2.150 18.635 2.260 ;
        RECT 17.945 1.285 18.850 1.515 ;
        RECT 20.805 1.230 21.035 2.260 ;
        RECT 10.410 0.770 12.235 1.000 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux4_4
MACRO gf180mcu_fd_sc_mcu9t5v0__nand2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.800 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.614500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.330 2.090 3.270 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.614500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 1.770 0.975 2.710 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.436200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 3.600 2.550 3.830 ;
        RECT 1.270 3.020 1.530 3.600 ;
        RECT 2.320 1.590 2.550 3.600 ;
        RECT 1.270 1.210 2.550 1.590 ;
        RECT 2.290 0.680 2.550 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 2.800 5.490 ;
        RECT 0.250 3.690 0.480 4.590 ;
        RECT 2.290 4.160 2.520 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 3.230 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 3.230 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 0.450 0.480 1.165 ;
        RECT 0.000 -0.450 2.800 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand2_1
MACRO gf180mcu_fd_sc_mcu9t5v0__nand2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.229000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.685 1.830 2.715 2.305 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.229000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.940 3.245 3.170 ;
        RECT 0.710 1.210 0.970 2.940 ;
        RECT 3.015 2.100 3.245 2.940 ;
        RECT 3.015 1.830 4.030 2.100 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.397200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 3.630 1.495 4.210 ;
        RECT 3.305 3.630 3.535 4.210 ;
        RECT 1.265 3.580 3.535 3.630 ;
        RECT 1.265 3.400 4.490 3.580 ;
        RECT 3.390 3.350 4.490 3.400 ;
        RECT 4.070 2.330 4.490 3.350 ;
        RECT 4.260 1.590 4.490 2.330 ;
        RECT 2.285 1.210 4.490 1.590 ;
        RECT 2.285 0.680 2.515 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.040 5.490 ;
        RECT 0.245 3.860 0.475 4.590 ;
        RECT 2.285 3.860 2.515 4.590 ;
        RECT 4.325 3.860 4.555 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 5.470 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 5.470 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.165 ;
        RECT 4.325 0.450 4.555 0.695 ;
        RECT 0.000 -0.450 5.040 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand2_2
MACRO gf180mcu_fd_sc_mcu9t5v0__nand2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.960 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.458000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.670 2.950 6.070 3.210 ;
        RECT 2.670 2.470 3.010 2.950 ;
        RECT 5.730 2.470 6.070 2.950 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.458000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.770 1.830 8.110 2.150 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.853800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 3.780 1.495 4.360 ;
        RECT 3.305 3.780 3.535 4.360 ;
        RECT 5.345 3.780 5.575 4.360 ;
        RECT 7.370 3.780 7.750 4.330 ;
        RECT 1.265 3.550 7.750 3.780 ;
        RECT 7.385 3.460 7.750 3.550 ;
        RECT 7.385 3.230 8.570 3.460 ;
        RECT 8.340 1.105 8.570 3.230 ;
        RECT 7.940 1.100 8.570 1.105 ;
        RECT 2.275 0.875 8.570 1.100 ;
        RECT 2.275 0.870 8.145 0.875 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 8.960 5.490 ;
        RECT 0.245 3.690 0.475 4.590 ;
        RECT 2.285 4.160 2.515 4.590 ;
        RECT 4.325 4.160 4.555 4.590 ;
        RECT 6.365 4.160 6.595 4.590 ;
        RECT 8.405 3.690 8.635 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.390 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.390 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.325 0.450 0.555 1.165 ;
        RECT 4.235 0.450 4.575 0.640 ;
        RECT 8.350 0.450 8.690 0.640 ;
        RECT 0.000 -0.450 8.960 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand2_4
MACRO gf180mcu_fd_sc_mcu9t5v0__nand3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 1.210 3.210 2.150 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.090 2.710 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.330 1.105 3.270 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.982400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 3.830 1.630 4.360 ;
        RECT 1.400 3.550 3.670 3.830 ;
        RECT 2.950 2.890 3.670 3.550 ;
        RECT 3.440 0.845 3.670 2.890 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 3.920 5.490 ;
        RECT 0.380 3.590 0.610 4.590 ;
        RECT 2.420 4.060 2.650 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.380 0.450 0.610 1.165 ;
        RECT 0.000 -0.450 3.920 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand3_1
MACRO gf180mcu_fd_sc_mcu9t5v0__nand3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.865 1.210 3.210 2.150 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.790 2.380 4.995 2.610 ;
        RECT 4.630 1.210 4.995 2.380 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.300 2.840 6.015 3.070 ;
        RECT 1.300 2.150 1.530 2.840 ;
        RECT 0.770 1.920 1.530 2.150 ;
        RECT 5.740 2.070 6.015 2.840 ;
        RECT 1.270 1.915 1.530 1.920 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.964000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 3.530 1.495 4.110 ;
        RECT 3.305 3.530 3.535 4.110 ;
        RECT 5.345 3.530 5.575 4.110 ;
        RECT 0.150 3.300 5.575 3.530 ;
        RECT 0.150 1.095 0.410 3.300 ;
        RECT 0.150 0.980 1.070 1.095 ;
        RECT 0.150 0.865 3.590 0.980 ;
        RECT 0.870 0.750 3.590 0.865 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.280 5.490 ;
        RECT 0.245 4.230 0.475 4.590 ;
        RECT 2.285 3.760 2.515 4.590 ;
        RECT 4.325 3.760 4.555 4.590 ;
        RECT 6.365 3.760 6.595 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.330 0.450 0.670 0.635 ;
        RECT 6.365 0.450 6.595 1.160 ;
        RECT 0.000 -0.450 7.280 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand3_2
MACRO gf180mcu_fd_sc_mcu9t5v0__nand3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.000 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.300 2.270 11.230 2.500 ;
        RECT 9.300 1.770 9.930 2.270 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.750 2.730 8.355 2.960 ;
        RECT 0.750 2.215 0.980 2.730 ;
        RECT 3.510 2.270 4.130 2.730 ;
        RECT 8.125 2.215 8.355 2.730 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.210 2.040 1.990 2.500 ;
        RECT 4.410 2.270 6.270 2.500 ;
        RECT 4.410 2.040 4.640 2.270 ;
        RECT 1.210 1.810 4.640 2.040 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.220000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 3.420 1.495 4.360 ;
        RECT 3.405 3.420 3.635 4.360 ;
        RECT 5.545 3.420 5.775 4.360 ;
        RECT 7.685 3.420 7.915 4.360 ;
        RECT 9.725 3.420 9.955 4.360 ;
        RECT 11.965 3.420 12.195 4.360 ;
        RECT 1.265 3.190 12.195 3.420 ;
        RECT 11.965 1.530 12.195 3.190 ;
        RECT 11.965 1.515 12.790 1.530 ;
        RECT 9.825 1.285 12.790 1.515 ;
        RECT 9.825 1.140 10.055 1.285 ;
        RECT 12.010 1.140 12.790 1.285 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.000 5.490 ;
        RECT 0.245 3.650 0.475 4.590 ;
        RECT 2.285 3.875 2.515 4.590 ;
        RECT 4.425 3.650 4.655 4.590 ;
        RECT 6.565 3.650 6.795 4.590 ;
        RECT 8.705 3.650 8.935 4.590 ;
        RECT 10.845 3.650 11.075 4.590 ;
        RECT 13.085 3.650 13.315 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.430 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.430 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.385 0.450 2.615 1.110 ;
        RECT 6.665 0.450 6.895 1.110 ;
        RECT 0.000 -0.450 14.000 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.350 3.075 1.580 ;
        RECT 0.245 0.770 0.475 1.350 ;
        RECT 2.845 1.000 3.075 1.350 ;
        RECT 4.525 1.350 9.170 1.580 ;
        RECT 4.525 1.000 4.755 1.350 ;
        RECT 2.845 0.770 4.755 1.000 ;
        RECT 8.940 0.910 9.170 1.350 ;
        RECT 10.890 0.910 11.230 1.055 ;
        RECT 13.185 0.910 13.415 1.580 ;
        RECT 8.940 0.680 13.415 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__nand3_4
MACRO gf180mcu_fd_sc_mcu9t5v0__nand4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.985 2.270 4.330 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.915 2.215 3.210 2.710 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.090 2.555 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 1.125 2.500 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.912000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.420 3.490 1.650 4.360 ;
        RECT 3.460 3.490 3.770 4.360 ;
        RECT 1.420 3.260 3.770 3.490 ;
        RECT 3.540 3.255 3.770 3.260 ;
        RECT 3.540 3.025 4.790 3.255 ;
        RECT 4.560 1.490 4.790 3.025 ;
        RECT 4.480 0.680 4.790 1.490 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.040 5.490 ;
        RECT 0.400 3.720 0.630 4.590 ;
        RECT 2.440 3.720 2.670 4.590 ;
        RECT 4.480 3.485 4.710 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 5.470 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 5.470 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 0.450 0.630 1.490 ;
        RECT 0.000 -0.450 5.040 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand4_1
MACRO gf180mcu_fd_sc_mcu9t5v0__nand4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.960 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 2.215 3.875 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.865 2.940 4.465 3.170 ;
        RECT 2.865 2.215 3.095 2.940 ;
        RECT 4.235 2.710 4.465 2.940 ;
        RECT 4.235 2.215 6.015 2.710 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.985 2.090 2.555 ;
        RECT 6.805 1.985 7.035 2.555 ;
        RECT 1.830 1.755 7.035 1.985 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.050 3.540 4.925 3.630 ;
        RECT 1.300 3.400 4.925 3.540 ;
        RECT 1.300 3.310 2.235 3.400 ;
        RECT 1.300 2.555 1.530 3.310 ;
        RECT 4.695 3.170 4.925 3.400 ;
        RECT 4.695 2.940 8.055 3.170 ;
        RECT 0.825 2.215 1.530 2.555 ;
        RECT 7.825 2.215 8.055 2.940 ;
        RECT 1.270 1.770 1.530 2.215 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.809600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 4.000 0.475 4.360 ;
        RECT 1.680 4.045 5.205 4.090 ;
        RECT 1.680 4.000 6.595 4.045 ;
        RECT 0.150 3.860 6.595 4.000 ;
        RECT 0.150 3.770 1.865 3.860 ;
        RECT 5.065 3.815 6.595 3.860 ;
        RECT 0.150 1.985 0.475 3.770 ;
        RECT 6.365 3.630 6.595 3.815 ;
        RECT 8.405 3.630 8.635 4.360 ;
        RECT 6.365 3.400 8.635 3.630 ;
        RECT 0.150 1.755 1.040 1.985 ;
        RECT 0.810 0.910 1.040 1.755 ;
        RECT 4.325 0.910 4.555 1.490 ;
        RECT 0.810 0.680 4.555 0.910 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 8.960 5.490 ;
        RECT 1.265 4.230 1.495 4.590 ;
        RECT 3.305 4.320 3.535 4.590 ;
        RECT 5.345 4.275 5.575 4.590 ;
        RECT 7.385 3.860 7.615 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.390 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.390 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 8.405 0.450 8.635 1.490 ;
        RECT 0.000 -0.450 8.960 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand4_2
MACRO gf180mcu_fd_sc_mcu9t5v0__nand4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.360 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.728000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.670 1.985 10.150 2.500 ;
        RECT 12.365 2.270 14.230 2.500 ;
        RECT 12.365 1.985 12.595 2.270 ;
        RECT 9.670 1.755 12.595 1.985 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.728000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.930 2.730 15.935 2.960 ;
        RECT 8.930 2.270 9.270 2.730 ;
        RECT 11.350 2.215 12.135 2.730 ;
        RECT 15.705 2.215 15.935 2.730 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.728000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.730 6.530 2.960 ;
        RECT 0.710 2.270 1.050 2.730 ;
        RECT 3.745 2.215 3.975 2.730 ;
        RECT 6.300 2.500 6.530 2.730 ;
        RECT 6.300 2.270 8.110 2.500 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.728000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.985 2.170 2.500 ;
        RECT 4.205 2.270 6.070 2.500 ;
        RECT 4.205 1.985 4.435 2.270 ;
        RECT 1.830 1.755 4.435 1.985 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.697600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 3.420 1.495 4.360 ;
        RECT 2.890 3.420 3.535 4.360 ;
        RECT 5.345 3.420 5.575 4.360 ;
        RECT 7.385 3.420 7.615 4.360 ;
        RECT 9.425 3.420 9.655 4.360 ;
        RECT 11.465 3.420 11.695 4.360 ;
        RECT 13.505 3.420 13.735 4.360 ;
        RECT 15.545 3.420 15.775 4.360 ;
        RECT 1.265 3.190 16.395 3.420 ;
        RECT 16.165 1.425 16.395 3.190 ;
        RECT 10.390 1.195 16.395 1.425 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.360 5.490 ;
        RECT 0.245 3.650 0.475 4.590 ;
        RECT 2.285 3.650 2.515 4.590 ;
        RECT 4.325 3.650 4.555 4.590 ;
        RECT 6.365 3.650 6.595 4.590 ;
        RECT 8.405 3.650 8.635 4.590 ;
        RECT 10.445 3.650 10.675 4.590 ;
        RECT 12.485 3.650 12.715 4.590 ;
        RECT 14.525 3.650 14.755 4.590 ;
        RECT 16.565 3.650 16.795 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 17.790 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 17.790 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.285 0.450 2.515 1.020 ;
        RECT 6.365 0.450 6.595 1.020 ;
        RECT 0.000 -0.450 17.360 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.260 10.160 1.490 ;
        RECT 0.245 0.680 0.475 1.260 ;
        RECT 4.325 0.680 4.555 1.260 ;
        RECT 9.930 0.965 10.160 1.260 ;
        RECT 9.930 0.735 16.850 0.965 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__nand4_4
MACRO gf180mcu_fd_sc_mcu9t5v0__nor2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.467000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.090 2.555 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.467000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.680 2.270 1.020 2.710 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.283600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.435 3.015 2.665 4.360 ;
        RECT 1.270 2.785 2.665 3.015 ;
        RECT 1.270 0.680 1.595 2.785 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 3.360 5.490 ;
        RECT 0.295 3.550 0.525 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 3.790 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 3.790 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.400 ;
        RECT 2.485 0.450 2.715 1.400 ;
        RECT 0.000 -0.450 3.360 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nor2_1
MACRO gf180mcu_fd_sc_mcu9t5v0__nor2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.934000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 2.270 2.140 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.934000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.875 2.940 3.950 3.170 ;
        RECT 0.875 2.215 1.105 2.940 ;
        RECT 3.510 2.270 3.950 2.940 ;
        RECT 3.510 1.770 3.770 2.270 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.999900 ;
    PORT
      LAYER Metal1 ;
        RECT 2.485 3.780 2.715 4.360 ;
        RECT 2.485 3.550 4.410 3.780 ;
        RECT 4.180 1.720 4.410 3.550 ;
        RECT 4.070 1.490 4.410 1.720 ;
        RECT 1.365 1.210 4.410 1.490 ;
        RECT 1.365 1.160 3.835 1.210 ;
        RECT 1.365 0.680 1.595 1.160 ;
        RECT 3.605 0.680 3.835 1.160 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.600 5.490 ;
        RECT 0.295 3.550 0.525 4.590 ;
        RECT 4.675 3.550 4.905 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.400 ;
        RECT 2.485 0.450 2.715 0.930 ;
        RECT 4.725 0.450 4.955 1.400 ;
        RECT 0.000 -0.450 5.600 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nor2_2
MACRO gf180mcu_fd_sc_mcu9t5v0__nor2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.868000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.060 2.270 3.810 2.500 ;
        RECT 3.580 2.000 3.810 2.270 ;
        RECT 4.630 2.270 6.620 2.500 ;
        RECT 4.630 2.000 4.890 2.270 ;
        RECT 3.580 1.770 4.890 2.000 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.868000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.600 2.730 7.080 2.960 ;
        RECT 2.600 2.500 2.830 2.730 ;
        RECT 1.200 2.270 2.830 2.500 ;
        RECT 4.040 2.270 4.380 2.730 ;
        RECT 6.850 2.500 7.080 2.730 ;
        RECT 6.850 2.270 8.860 2.500 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.091300 ;
    PORT
      LAYER Metal1 ;
        RECT 2.485 3.420 2.715 4.360 ;
        RECT 6.915 3.420 7.145 4.360 ;
        RECT 0.710 3.190 7.145 3.420 ;
        RECT 0.710 1.490 0.970 3.190 ;
        RECT 0.710 1.260 8.315 1.490 ;
        RECT 1.365 0.680 1.595 1.260 ;
        RECT 3.605 0.680 3.835 1.260 ;
        RECT 5.845 0.680 6.075 1.260 ;
        RECT 8.085 0.680 8.315 1.260 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 10.080 5.490 ;
        RECT 0.295 3.650 0.525 4.590 ;
        RECT 4.675 3.650 4.905 4.590 ;
        RECT 9.155 3.650 9.385 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 10.510 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.020 ;
        RECT 4.725 0.450 4.955 1.020 ;
        RECT 6.965 0.450 7.195 1.020 ;
        RECT 9.205 0.450 9.435 1.400 ;
        RECT 0.000 -0.450 10.080 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nor2_4
MACRO gf180mcu_fd_sc_mcu9t5v0__nor3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 1.770 3.210 2.555 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 2.270 2.140 2.710 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.215 1.015 2.710 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.563600 ;
    PORT
      LAYER Metal1 ;
        RECT 3.505 1.480 3.835 4.360 ;
        RECT 1.365 1.250 3.835 1.480 ;
        RECT 1.365 0.680 1.595 1.250 ;
        RECT 3.605 0.680 3.835 1.250 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 4.480 5.490 ;
        RECT 0.345 3.550 0.575 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.020 ;
        RECT 2.485 0.450 2.715 1.020 ;
        RECT 0.000 -0.450 4.480 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nor3_1
MACRO gf180mcu_fd_sc_mcu9t5v0__nor3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.475 2.215 3.770 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.940 5.445 3.170 ;
        RECT 1.830 2.215 2.135 2.940 ;
        RECT 5.215 2.215 5.445 2.940 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 3.400 6.570 3.630 ;
        RECT 1.265 2.215 1.495 3.400 ;
        RECT 6.310 2.215 6.570 3.400 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.651400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.805 3.930 3.840 4.160 ;
        RECT 0.805 1.590 1.035 3.930 ;
        RECT 0.245 1.480 1.035 1.590 ;
        RECT 0.245 1.250 7.195 1.480 ;
        RECT 0.245 1.210 2.715 1.250 ;
        RECT 0.245 0.680 0.475 1.210 ;
        RECT 2.485 0.680 2.715 1.210 ;
        RECT 4.725 0.680 4.955 1.250 ;
        RECT 6.965 0.680 7.195 1.250 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.840 5.490 ;
        RECT 0.345 3.875 0.575 4.590 ;
        RECT 6.865 3.875 7.095 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 8.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.980 ;
        RECT 3.605 0.450 3.835 1.020 ;
        RECT 5.845 0.450 6.075 1.020 ;
        RECT 0.000 -0.450 7.840 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nor3_2
MACRO gf180mcu_fd_sc_mcu9t5v0__nor3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.800 1.710 11.730 2.150 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.825 2.895 6.975 3.125 ;
        RECT 0.825 2.325 1.055 2.895 ;
        RECT 3.510 2.380 4.330 2.895 ;
        RECT 6.745 2.610 6.975 2.895 ;
        RECT 6.745 2.380 8.810 2.610 ;
        RECT 3.510 2.330 3.770 2.380 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.940 2.000 3.280 2.610 ;
        RECT 6.285 2.150 6.515 2.665 ;
        RECT 4.070 2.000 6.515 2.150 ;
        RECT 2.940 1.770 6.515 2.000 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.734000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.325 2.880 10.555 3.900 ;
        RECT 11.910 3.090 12.695 3.900 ;
        RECT 11.910 2.880 12.190 3.090 ;
        RECT 10.325 2.650 12.190 2.880 ;
        RECT 11.960 1.480 12.190 2.650 ;
        RECT 1.365 1.250 12.795 1.480 ;
        RECT 1.365 0.680 1.595 1.250 ;
        RECT 3.605 0.680 3.835 1.250 ;
        RECT 5.845 0.680 6.075 1.250 ;
        RECT 8.085 0.680 8.315 1.250 ;
        RECT 10.325 0.680 10.555 1.250 ;
        RECT 12.565 0.680 12.795 1.250 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.560 5.490 ;
        RECT 2.385 3.825 2.615 4.590 ;
        RECT 6.865 3.815 7.095 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.020 ;
        RECT 2.485 0.450 2.715 1.020 ;
        RECT 4.725 0.450 4.955 1.020 ;
        RECT 6.965 0.450 7.195 1.020 ;
        RECT 9.205 0.450 9.435 1.020 ;
        RECT 11.445 0.450 11.675 1.020 ;
        RECT 13.685 0.450 13.915 1.020 ;
        RECT 0.000 -0.450 14.560 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.585 0.475 3.920 ;
        RECT 4.625 3.585 4.855 4.165 ;
        RECT 7.375 4.130 13.815 4.360 ;
        RECT 7.375 3.585 7.605 4.130 ;
        RECT 0.245 3.355 7.605 3.585 ;
        RECT 0.245 3.110 0.475 3.355 ;
        RECT 11.345 3.110 11.575 4.130 ;
        RECT 13.585 3.110 13.815 4.130 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__nor3_4
MACRO gf180mcu_fd_sc_mcu9t5v0__nor4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.311000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.070 1.770 4.330 2.555 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.311000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.920 2.270 3.260 2.710 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.311000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 2.270 2.140 2.710 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.311000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.215 1.015 2.710 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.491600 ;
    PORT
      LAYER Metal1 ;
        RECT 4.625 3.015 4.855 4.360 ;
        RECT 3.510 2.785 4.855 3.015 ;
        RECT 3.510 1.440 3.835 2.785 ;
        RECT 1.365 1.210 3.835 1.440 ;
        RECT 1.365 0.680 1.595 1.210 ;
        RECT 3.605 0.680 3.835 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.600 5.490 ;
        RECT 0.345 3.550 0.575 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.005 ;
        RECT 2.485 0.450 2.715 0.980 ;
        RECT 4.725 0.450 4.955 1.005 ;
        RECT 0.000 -0.450 5.600 0.450 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nor4_1
MACRO gf180mcu_fd_sc_mcu9t5v0__nor4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.622000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.870 2.150 7.130 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.622000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.340 2.940 9.120 3.170 ;
        RECT 6.340 2.555 6.570 2.940 ;
        RECT 5.770 1.770 6.570 2.555 ;
        RECT 8.890 2.215 9.120 2.940 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.622000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.930 2.785 4.510 3.015 ;
        RECT 0.930 2.215 1.160 2.785 ;
        RECT 4.070 1.770 4.510 2.785 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.622000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.090 2.555 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.718200 ;
    PORT
      LAYER Metal1 ;
        RECT 7.280 3.630 7.510 3.890 ;
        RECT 5.190 3.400 7.510 3.630 ;
        RECT 5.190 1.455 5.450 3.400 ;
        RECT 1.370 1.225 8.680 1.455 ;
        RECT 1.370 0.680 1.600 1.225 ;
        RECT 3.610 1.210 6.440 1.225 ;
        RECT 3.610 0.680 3.840 1.210 ;
        RECT 6.210 0.680 6.440 1.210 ;
        RECT 8.450 0.680 8.680 1.225 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 10.080 5.490 ;
        RECT 2.440 3.705 2.670 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 10.510 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 0.450 0.480 1.020 ;
        RECT 2.490 0.450 2.720 0.995 ;
        RECT 4.910 0.450 5.140 0.980 ;
        RECT 7.330 0.450 7.560 0.995 ;
        RECT 9.570 0.450 9.800 0.995 ;
        RECT 0.000 -0.450 10.080 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.350 4.130 2.210 4.360 ;
        RECT 0.350 3.550 0.580 4.130 ;
        RECT 1.980 3.475 2.210 4.130 ;
        RECT 2.900 4.130 9.700 4.360 ;
        RECT 2.900 3.475 3.130 4.130 ;
        RECT 9.470 3.550 9.700 4.130 ;
        RECT 1.980 3.245 3.130 3.475 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__nor4_2
MACRO gf180mcu_fd_sc_mcu9t5v0__nor4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.244000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.465 2.215 17.460 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.244000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.870 1.985 11.100 2.555 ;
        RECT 19.550 1.985 20.010 2.555 ;
        RECT 10.870 1.755 20.010 1.985 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.244000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 2.785 7.700 3.015 ;
        RECT 1.100 2.150 1.330 2.785 ;
        RECT 4.590 2.215 4.820 2.785 ;
        RECT 7.470 2.500 7.700 2.785 ;
        RECT 7.470 2.270 9.715 2.500 ;
        RECT 0.710 1.770 1.330 2.150 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.244000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.480 1.985 3.710 2.555 ;
        RECT 6.780 1.985 7.240 2.555 ;
        RECT 3.480 1.755 7.240 1.985 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.389400 ;
    PORT
      LAYER Metal1 ;
        RECT 12.890 3.320 13.120 3.900 ;
        RECT 17.810 3.320 18.040 3.900 ;
        RECT 12.890 3.090 20.635 3.320 ;
        RECT 20.405 1.590 20.635 3.090 ;
        RECT 20.175 1.455 20.635 1.590 ;
        RECT 1.680 1.225 5.910 1.455 ;
        RECT 1.680 0.680 1.910 1.225 ;
        RECT 3.920 0.680 4.150 1.225 ;
        RECT 5.680 0.910 5.910 1.225 ;
        RECT 6.520 1.225 20.635 1.455 ;
        RECT 6.520 0.910 6.750 1.225 ;
        RECT 5.680 0.680 6.750 0.910 ;
        RECT 8.760 0.680 8.990 1.225 ;
        RECT 11.360 0.680 11.590 1.225 ;
        RECT 13.960 0.680 14.190 1.225 ;
        RECT 16.560 0.680 16.790 1.225 ;
        RECT 19.160 1.210 20.635 1.225 ;
        RECT 19.160 0.680 19.390 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 21.280 5.490 ;
        RECT 2.750 3.705 2.980 4.590 ;
        RECT 7.590 3.705 7.820 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 21.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.560 0.450 0.790 0.995 ;
        RECT 2.800 0.450 3.030 0.995 ;
        RECT 5.220 0.450 5.450 0.995 ;
        RECT 7.640 0.450 7.870 0.995 ;
        RECT 10.060 0.450 10.290 0.995 ;
        RECT 12.660 0.450 12.890 0.995 ;
        RECT 15.260 0.450 15.490 0.970 ;
        RECT 17.860 0.450 18.090 0.995 ;
        RECT 20.460 0.450 20.690 0.980 ;
        RECT 0.000 -0.450 21.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.660 4.130 2.520 4.360 ;
        RECT 0.660 3.550 0.890 4.130 ;
        RECT 2.290 3.475 2.520 4.130 ;
        RECT 5.170 3.475 5.400 4.360 ;
        RECT 8.050 4.130 20.590 4.360 ;
        RECT 8.050 3.475 8.280 4.130 ;
        RECT 15.210 3.550 15.440 4.130 ;
        RECT 20.360 3.550 20.590 4.130 ;
        RECT 2.290 3.245 8.280 3.475 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__nor4_4
MACRO gf180mcu_fd_sc_mcu9t5v0__oai21_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai21_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.090 2.555 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.680 2.270 1.020 2.710 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.614500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 2.270 3.290 2.710 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.911900 ;
    PORT
      LAYER Metal1 ;
        RECT 2.385 3.015 2.615 4.360 ;
        RECT 1.270 2.785 2.615 3.015 ;
        RECT 1.270 1.140 1.595 2.785 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 4.480 5.490 ;
        RECT 0.295 3.550 0.525 4.590 ;
        RECT 3.585 3.550 3.815 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.605 0.450 3.835 1.655 ;
        RECT 0.000 -0.450 4.480 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 0.910 0.475 1.655 ;
        RECT 2.485 0.910 2.715 1.655 ;
        RECT 0.245 0.680 2.715 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai21_1
MACRO gf180mcu_fd_sc_mcu9t5v0__oai21_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai21_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.035 2.215 4.330 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 2.940 6.515 3.170 ;
        RECT 2.950 2.270 3.310 2.940 ;
        RECT 6.285 2.215 6.515 2.940 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.229000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 2.270 1.070 2.650 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.362800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.630 1.595 4.320 ;
        RECT 4.675 3.630 4.905 4.360 ;
        RECT 1.365 3.400 6.975 3.630 ;
        RECT 6.745 1.950 6.975 3.400 ;
        RECT 3.605 1.720 6.975 1.950 ;
        RECT 3.605 1.140 3.835 1.720 ;
        RECT 5.190 1.140 6.075 1.720 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.840 5.490 ;
        RECT 0.345 3.665 0.575 4.590 ;
        RECT 2.385 3.860 2.615 4.590 ;
        RECT 6.865 3.860 7.095 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 8.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.490 ;
        RECT 0.000 -0.450 7.840 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.720 2.715 1.950 ;
        RECT 0.245 0.680 0.475 1.720 ;
        RECT 2.485 0.910 2.715 1.720 ;
        RECT 4.725 0.910 4.955 1.490 ;
        RECT 6.965 0.910 7.195 1.490 ;
        RECT 2.485 0.680 7.195 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai21_2
MACRO gf180mcu_fd_sc_mcu9t5v0__oai21_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai21_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.060 2.270 3.770 2.500 ;
        RECT 3.510 2.040 3.770 2.270 ;
        RECT 4.610 2.270 6.570 2.500 ;
        RECT 4.610 2.040 4.840 2.270 ;
        RECT 3.510 1.810 4.840 2.040 ;
        RECT 3.510 1.770 3.770 1.810 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.600 2.730 7.030 2.960 ;
        RECT 2.600 2.500 2.830 2.730 ;
        RECT 1.250 2.270 2.830 2.500 ;
        RECT 4.040 2.270 4.380 2.730 ;
        RECT 6.800 2.500 7.030 2.730 ;
        RECT 6.800 2.270 8.810 2.500 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.458000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.270 2.270 12.850 2.500 ;
        RECT 11.350 1.770 11.610 2.270 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.798600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.485 3.420 2.715 4.360 ;
        RECT 6.915 3.420 7.145 4.360 ;
        RECT 10.325 3.420 10.555 4.360 ;
        RECT 12.515 3.420 12.745 4.360 ;
        RECT 0.790 3.190 12.745 3.420 ;
        RECT 0.790 2.040 1.020 3.190 ;
        RECT 0.790 1.810 3.210 2.040 ;
        RECT 1.365 1.140 1.595 1.810 ;
        RECT 2.950 1.480 3.210 1.810 ;
        RECT 3.935 1.480 8.315 1.570 ;
        RECT 2.950 1.340 8.315 1.480 ;
        RECT 2.950 1.140 4.120 1.340 ;
        RECT 5.845 1.140 6.075 1.340 ;
        RECT 8.085 1.140 8.315 1.340 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.560 5.490 ;
        RECT 0.345 3.650 0.575 4.590 ;
        RECT 4.675 3.650 4.905 4.590 ;
        RECT 9.105 3.650 9.335 4.590 ;
        RECT 11.345 3.650 11.575 4.590 ;
        RECT 13.635 3.650 13.865 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 10.325 0.450 10.555 1.195 ;
        RECT 12.565 0.450 12.795 1.110 ;
        RECT 0.000 -0.450 14.560 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 0.910 0.475 1.580 ;
        RECT 2.485 0.910 2.715 1.580 ;
        RECT 9.205 1.540 11.150 1.655 ;
        RECT 11.775 1.540 13.915 1.580 ;
        RECT 9.205 1.425 13.915 1.540 ;
        RECT 4.725 0.910 4.955 1.110 ;
        RECT 6.965 0.910 7.195 1.110 ;
        RECT 9.205 0.910 9.435 1.425 ;
        RECT 10.950 1.350 13.915 1.425 ;
        RECT 10.950 1.310 11.905 1.350 ;
        RECT 0.245 0.680 9.435 0.910 ;
        RECT 11.445 0.730 11.905 1.310 ;
        RECT 13.685 0.770 13.915 1.350 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai21_4
MACRO gf180mcu_fd_sc_mcu9t5v0__oai22_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai22_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 1.770 3.210 2.555 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.070 1.770 4.330 2.555 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 2.270 2.140 2.710 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.215 1.015 3.270 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.535 3.015 2.765 4.360 ;
        RECT 2.535 2.785 3.835 3.015 ;
        RECT 3.510 1.140 3.835 2.785 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.600 5.490 ;
        RECT 0.345 3.550 0.575 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.525 ;
        RECT 0.000 -0.450 5.600 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.755 2.715 1.985 ;
        RECT 0.245 0.715 0.475 1.755 ;
        RECT 2.485 0.910 2.715 1.755 ;
        RECT 4.725 0.910 4.955 1.525 ;
        RECT 2.485 0.680 4.955 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai22_1
MACRO gf180mcu_fd_sc_mcu9t5v0__oai22_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai22_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.280 2.270 6.620 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.350 2.940 8.755 3.170 ;
        RECT 5.350 2.270 5.690 2.940 ;
        RECT 6.870 2.215 8.755 2.940 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.750 2.270 2.090 2.710 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.870 2.940 4.330 3.170 ;
        RECT 0.870 2.270 1.210 2.940 ;
        RECT 2.390 2.270 4.330 2.940 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.733500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.535 3.630 2.765 4.360 ;
        RECT 6.915 3.630 7.145 4.360 ;
        RECT 2.535 3.400 9.215 3.630 ;
        RECT 8.985 1.985 9.215 3.400 ;
        RECT 5.845 1.755 9.215 1.985 ;
        RECT 5.845 1.140 6.075 1.755 ;
        RECT 7.990 1.140 8.315 1.755 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 10.080 5.490 ;
        RECT 0.345 3.860 0.575 4.590 ;
        RECT 4.625 3.860 4.855 4.590 ;
        RECT 9.105 3.860 9.335 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 10.510 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.525 ;
        RECT 3.605 0.450 3.835 1.055 ;
        RECT 0.000 -0.450 10.080 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.755 4.955 1.985 ;
        RECT 0.245 0.715 0.475 1.755 ;
        RECT 2.485 1.285 4.955 1.755 ;
        RECT 4.725 0.910 4.955 1.285 ;
        RECT 6.965 0.910 7.195 1.525 ;
        RECT 9.205 0.910 9.435 1.525 ;
        RECT 4.725 0.680 9.435 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai22_2
MACRO gf180mcu_fd_sc_mcu9t5v0__oai22_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai22_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.730 1.985 11.340 2.500 ;
        RECT 13.515 2.270 15.530 2.500 ;
        RECT 13.515 1.985 13.745 2.270 ;
        RECT 10.730 1.755 13.745 1.985 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.885 2.730 17.715 2.960 ;
        RECT 9.885 2.215 10.115 2.730 ;
        RECT 12.470 2.215 13.285 2.730 ;
        RECT 17.485 2.215 17.715 2.730 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.110 2.040 3.450 2.500 ;
        RECT 4.810 2.270 6.570 2.500 ;
        RECT 4.810 2.150 5.040 2.270 ;
        RECT 4.580 2.040 5.040 2.150 ;
        RECT 3.110 1.770 5.040 2.040 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.875 2.730 7.030 2.960 ;
        RECT 0.875 2.215 1.105 2.730 ;
        RECT 4.040 2.270 4.380 2.730 ;
        RECT 6.800 2.500 7.030 2.730 ;
        RECT 6.800 2.270 8.810 2.500 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.558500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.585 3.420 2.815 4.360 ;
        RECT 6.865 3.420 7.095 4.360 ;
        RECT 11.395 3.420 11.625 4.360 ;
        RECT 15.975 3.830 16.205 4.360 ;
        RECT 15.975 3.450 18.330 3.830 ;
        RECT 15.975 3.420 18.175 3.450 ;
        RECT 2.585 3.190 18.175 3.420 ;
        RECT 17.945 1.475 18.175 3.190 ;
        RECT 10.270 1.245 18.175 1.475 ;
        RECT 10.270 1.140 10.610 1.245 ;
        RECT 12.510 1.140 15.090 1.245 ;
        RECT 16.990 1.140 18.175 1.245 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 19.040 5.490 ;
        RECT 0.295 3.550 0.525 4.590 ;
        RECT 4.675 3.650 4.905 4.590 ;
        RECT 9.105 3.650 9.335 4.590 ;
        RECT 13.635 3.650 13.865 4.590 ;
        RECT 18.065 4.060 18.295 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 19.470 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 19.470 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.070 ;
        RECT 3.605 0.450 3.835 1.070 ;
        RECT 5.845 0.450 6.075 1.070 ;
        RECT 8.085 0.450 8.315 1.070 ;
        RECT 0.000 -0.450 19.040 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.310 9.435 1.540 ;
        RECT 0.245 0.730 0.475 1.310 ;
        RECT 2.485 0.730 2.715 1.310 ;
        RECT 4.725 0.730 4.955 1.310 ;
        RECT 6.965 0.730 7.195 1.310 ;
        RECT 9.205 0.910 9.435 1.310 ;
        RECT 11.390 0.910 11.730 1.015 ;
        RECT 15.870 0.910 16.210 1.015 ;
        RECT 18.405 0.910 18.635 1.540 ;
        RECT 9.205 0.680 18.635 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai22_4
MACRO gf180mcu_fd_sc_mcu9t5v0__oai31_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai31_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.135 2.555 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.920 1.770 3.260 2.500 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.990 1.770 4.330 2.500 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.614500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 1.770 0.970 2.500 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.525600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.465 3.830 1.695 4.360 ;
        RECT 1.465 3.450 2.650 3.830 ;
        RECT 2.420 1.540 2.650 3.450 ;
        RECT 2.420 1.310 4.955 1.540 ;
        RECT 2.420 1.140 2.770 1.310 ;
        RECT 4.725 0.730 4.955 1.310 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.600 5.490 ;
        RECT 0.245 3.550 0.475 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.540 ;
        RECT 0.000 -0.450 5.600 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 0.910 1.595 1.540 ;
        RECT 3.605 0.910 3.835 1.070 ;
        RECT 1.365 0.680 3.835 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai31_1
MACRO gf180mcu_fd_sc_mcu9t5v0__oai31_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai31_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.630 2.270 5.500 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.040 2.150 4.380 2.500 ;
        RECT 3.510 2.040 4.380 2.150 ;
        RECT 6.045 2.215 7.685 2.555 ;
        RECT 6.045 2.040 6.275 2.215 ;
        RECT 3.510 1.810 6.275 2.040 ;
        RECT 3.510 1.770 3.770 1.810 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.055 2.940 8.220 3.170 ;
        RECT 3.055 2.215 3.285 2.940 ;
        RECT 7.990 2.710 8.220 2.940 ;
        RECT 7.990 2.215 8.755 2.710 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.229000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.675 2.215 0.970 2.710 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.131450 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.630 1.595 4.360 ;
        RECT 5.795 3.630 6.025 4.360 ;
        RECT 1.365 3.400 9.215 3.630 ;
        RECT 8.985 1.935 9.215 3.400 ;
        RECT 6.505 1.705 9.215 1.935 ;
        RECT 6.505 1.580 6.735 1.705 ;
        RECT 3.935 1.540 6.735 1.580 ;
        RECT 3.605 1.350 6.735 1.540 ;
        RECT 3.605 1.140 4.065 1.350 ;
        RECT 5.845 1.140 6.735 1.350 ;
        RECT 7.430 1.140 8.315 1.705 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 10.080 5.490 ;
        RECT 0.295 3.860 0.525 4.590 ;
        RECT 2.385 3.860 2.615 4.590 ;
        RECT 9.105 3.860 9.335 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 10.510 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.525 ;
        RECT 0.000 -0.450 10.080 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.755 2.715 1.985 ;
        RECT 0.245 0.845 0.475 1.755 ;
        RECT 2.485 0.910 2.715 1.755 ;
        RECT 4.725 0.910 4.955 1.120 ;
        RECT 6.965 0.910 7.195 1.185 ;
        RECT 9.440 0.910 9.670 1.655 ;
        RECT 2.485 0.680 9.670 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai31_2
MACRO gf180mcu_fd_sc_mcu9t5v0__oai31_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai31_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.590 2.270 8.250 2.500 ;
        RECT 7.990 2.000 8.250 2.270 ;
        RECT 10.160 2.270 11.100 2.500 ;
        RECT 10.160 2.000 10.390 2.270 ;
        RECT 7.990 1.770 10.390 2.000 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.355 2.730 13.235 2.960 ;
        RECT 5.355 2.215 5.585 2.730 ;
        RECT 9.590 2.270 9.930 2.730 ;
        RECT 13.005 2.215 13.235 2.730 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 2.270 3.890 2.500 ;
        RECT 1.270 1.770 1.530 2.270 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.458000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.270 2.270 17.850 2.710 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 8.509650 ;
    PORT
      LAYER Metal1 ;
        RECT 6.960 3.605 11.625 3.890 ;
        RECT 11.395 3.420 11.625 3.605 ;
        RECT 15.325 3.420 15.555 4.360 ;
        RECT 11.395 3.320 15.555 3.420 ;
        RECT 17.515 3.320 17.745 4.360 ;
        RECT 11.395 3.190 17.745 3.320 ;
        RECT 13.465 3.090 17.745 3.190 ;
        RECT 13.465 1.985 13.695 3.090 ;
        RECT 10.620 1.755 13.695 1.985 ;
        RECT 1.695 1.540 7.825 1.605 ;
        RECT 10.620 1.540 10.850 1.755 ;
        RECT 1.365 1.375 10.850 1.540 ;
        RECT 1.365 1.140 1.860 1.375 ;
        RECT 3.550 1.140 3.890 1.375 ;
        RECT 5.190 1.140 6.130 1.375 ;
        RECT 7.660 1.310 10.850 1.375 ;
        RECT 7.660 1.140 8.370 1.310 ;
        RECT 10.270 1.140 10.850 1.310 ;
        RECT 12.565 1.140 12.795 1.755 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 19.600 5.490 ;
        RECT 1.365 3.550 1.595 4.590 ;
        RECT 3.555 3.550 3.785 4.590 ;
        RECT 14.305 3.875 14.535 4.590 ;
        RECT 16.495 3.550 16.725 4.590 ;
        RECT 18.635 3.550 18.865 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 20.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 20.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 15.325 0.450 15.555 1.580 ;
        RECT 17.565 0.450 17.795 1.580 ;
        RECT 0.000 -0.450 19.600 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.320 0.575 4.360 ;
        RECT 2.485 3.320 2.715 4.360 ;
        RECT 4.935 4.120 13.870 4.350 ;
        RECT 4.935 3.320 5.165 4.120 ;
        RECT 0.345 3.090 5.165 3.320 ;
        RECT 13.925 1.810 18.915 2.040 ;
        RECT 0.245 0.910 0.475 1.615 ;
        RECT 2.485 0.910 2.715 1.145 ;
        RECT 4.725 0.910 4.955 1.145 ;
        RECT 6.965 0.910 7.195 1.145 ;
        RECT 9.150 0.910 9.490 1.080 ;
        RECT 11.445 0.910 11.675 1.525 ;
        RECT 13.925 0.910 14.155 1.810 ;
        RECT 0.245 0.680 14.155 0.910 ;
        RECT 16.445 0.805 16.675 1.810 ;
        RECT 18.685 0.805 18.915 1.810 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai31_4
MACRO gf180mcu_fd_sc_mcu9t5v0__oai32_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai32_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.920 2.270 3.260 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 2.270 2.140 2.710 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.215 1.015 2.710 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.070 1.770 4.330 2.555 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.190 1.770 5.450 2.555 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.655 3.015 3.885 4.360 ;
        RECT 3.655 2.785 4.955 3.015 ;
        RECT 4.630 1.140 4.955 2.785 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 6.720 5.490 ;
        RECT 0.345 3.550 0.575 4.590 ;
        RECT 5.745 3.550 5.975 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.150 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.150 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.580 ;
        RECT 2.485 0.450 2.715 1.580 ;
        RECT 0.000 -0.450 6.720 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 1.810 3.835 2.040 ;
        RECT 1.365 0.770 1.595 1.810 ;
        RECT 3.605 0.910 3.835 1.810 ;
        RECT 5.845 0.910 6.075 1.580 ;
        RECT 3.605 0.680 6.075 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai32_1
MACRO gf180mcu_fd_sc_mcu9t5v0__oai32_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai32_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.320 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.920 2.270 3.260 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.940 2.270 2.690 2.500 ;
        RECT 2.460 2.040 2.690 2.270 ;
        RECT 4.630 2.270 5.450 2.500 ;
        RECT 4.630 2.040 4.890 2.270 ;
        RECT 2.460 1.810 4.890 2.040 ;
        RECT 4.630 1.770 4.890 1.810 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.940 5.910 3.170 ;
        RECT 0.710 2.215 1.015 2.940 ;
        RECT 5.680 2.500 5.910 2.940 ;
        RECT 5.680 2.270 6.570 2.500 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.515 2.215 8.810 2.710 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.430 2.940 10.995 3.170 ;
        RECT 7.430 2.215 7.735 2.940 ;
        RECT 10.765 2.215 10.995 2.940 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.655 3.645 3.885 4.355 ;
        RECT 9.155 3.645 9.385 4.340 ;
        RECT 3.655 3.415 11.455 3.645 ;
        RECT 11.225 1.985 11.455 3.415 ;
        RECT 7.990 1.755 11.455 1.985 ;
        RECT 7.990 1.140 8.315 1.755 ;
        RECT 10.325 1.140 10.555 1.755 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 12.320 5.490 ;
        RECT 0.345 3.875 0.575 4.590 ;
        RECT 6.865 3.875 7.095 4.590 ;
        RECT 11.345 3.875 11.575 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 12.750 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.750 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.095 ;
        RECT 3.605 0.450 3.835 1.095 ;
        RECT 5.845 0.450 6.075 1.095 ;
        RECT 0.000 -0.450 12.320 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.540 4.475 1.565 ;
        RECT 5.055 1.540 7.195 1.565 ;
        RECT 0.245 1.335 7.195 1.540 ;
        RECT 0.245 0.755 0.475 1.335 ;
        RECT 2.485 0.755 2.715 1.335 ;
        RECT 4.370 1.310 5.160 1.335 ;
        RECT 4.725 0.730 5.160 1.310 ;
        RECT 6.965 0.910 7.195 1.335 ;
        RECT 9.205 0.910 9.435 1.525 ;
        RECT 11.685 0.910 11.915 1.565 ;
        RECT 6.965 0.680 11.915 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai32_2
MACRO gf180mcu_fd_sc_mcu9t5v0__oai32_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai32_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.080 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.670 2.270 13.055 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.080 2.785 4.475 3.015 ;
        RECT 1.080 2.215 1.310 2.785 ;
        RECT 4.245 2.500 4.475 2.785 ;
        RECT 6.870 2.785 9.010 3.015 ;
        RECT 6.870 2.500 7.130 2.785 ;
        RECT 4.245 2.270 7.130 2.500 ;
        RECT 8.780 2.215 9.010 2.785 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.370 2.040 3.600 2.555 ;
        RECT 7.430 2.040 7.690 2.555 ;
        RECT 3.370 1.810 7.690 2.040 ;
        RECT 7.430 1.770 7.690 1.810 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 17.275 2.040 17.615 2.500 ;
        RECT 20.310 2.270 20.785 2.500 ;
        RECT 20.310 2.040 20.570 2.270 ;
        RECT 17.275 1.810 20.570 2.040 ;
        RECT 20.310 1.770 20.570 1.810 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 18.630 2.960 18.890 3.270 ;
        RECT 15.305 2.730 18.075 2.960 ;
        RECT 15.305 2.500 15.535 2.730 ;
        RECT 15.035 2.270 15.535 2.500 ;
        RECT 17.845 2.500 18.075 2.730 ;
        RECT 18.630 2.730 22.590 2.960 ;
        RECT 18.630 2.500 18.860 2.730 ;
        RECT 17.845 2.270 18.860 2.500 ;
        RECT 22.360 2.215 22.590 2.730 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.467000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.530 3.320 10.760 3.900 ;
        RECT 12.570 3.320 12.800 3.900 ;
        RECT 16.700 3.770 21.310 4.000 ;
        RECT 16.700 3.450 17.210 3.770 ;
        RECT 16.700 3.420 16.930 3.450 ;
        RECT 14.925 3.320 16.930 3.420 ;
        RECT 10.530 3.190 16.930 3.320 ;
        RECT 21.080 3.420 21.310 3.770 ;
        RECT 21.080 3.190 23.050 3.420 ;
        RECT 10.530 3.090 15.115 3.190 ;
        RECT 15.530 1.540 20.070 1.570 ;
        RECT 22.820 1.565 23.050 3.190 ;
        RECT 20.675 1.540 23.050 1.565 ;
        RECT 15.530 1.340 23.050 1.540 ;
        RECT 15.530 1.140 15.760 1.340 ;
        RECT 17.770 1.140 18.000 1.340 ;
        RECT 19.955 1.335 23.050 1.340 ;
        RECT 19.955 1.140 20.780 1.335 ;
        RECT 22.250 1.140 23.050 1.335 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 24.080 5.490 ;
        RECT 2.590 3.705 2.820 4.590 ;
        RECT 7.070 3.705 7.300 4.590 ;
        RECT 14.510 3.560 14.740 4.590 ;
        RECT 18.840 4.345 19.070 4.590 ;
        RECT 23.280 3.090 23.510 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 24.510 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 24.510 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.570 0.450 1.800 1.110 ;
        RECT 3.810 0.450 4.040 1.110 ;
        RECT 6.050 0.450 6.280 1.110 ;
        RECT 8.290 0.450 8.520 1.110 ;
        RECT 10.530 0.450 10.760 1.110 ;
        RECT 12.770 0.450 13.000 1.110 ;
        RECT 0.000 -0.450 24.080 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 7.530 4.130 14.020 4.360 ;
        RECT 0.500 3.475 0.730 3.900 ;
        RECT 4.880 3.475 5.110 3.900 ;
        RECT 7.530 3.475 7.760 4.130 ;
        RECT 11.550 3.550 11.780 4.130 ;
        RECT 13.790 3.550 14.020 4.130 ;
        RECT 0.500 3.245 7.760 3.475 ;
        RECT 0.500 3.090 0.730 3.245 ;
        RECT 4.880 3.090 5.110 3.245 ;
        RECT 0.450 1.540 7.300 1.580 ;
        RECT 7.820 1.540 14.120 1.580 ;
        RECT 0.450 1.350 14.120 1.540 ;
        RECT 0.450 0.770 0.680 1.350 ;
        RECT 2.690 0.770 2.920 1.350 ;
        RECT 4.930 0.770 5.160 1.350 ;
        RECT 7.170 1.310 7.950 1.350 ;
        RECT 7.170 0.730 7.400 1.310 ;
        RECT 9.410 0.770 9.640 1.350 ;
        RECT 11.650 0.770 11.880 1.350 ;
        RECT 13.890 0.910 14.120 1.350 ;
        RECT 16.650 0.910 16.880 1.110 ;
        RECT 18.890 0.910 19.120 1.110 ;
        RECT 21.130 0.910 21.360 1.105 ;
        RECT 23.370 0.910 23.600 1.580 ;
        RECT 13.890 0.680 23.600 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai32_4
MACRO gf180mcu_fd_sc_mcu9t5v0__oai33_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai33_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.070 1.770 4.330 2.555 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.190 2.215 5.450 3.270 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.230 2.270 6.570 2.710 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.920 2.270 3.260 2.710 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 2.270 2.140 2.710 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.215 1.015 2.710 ;
    END
  END B3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.401800 ;
    PORT
      LAYER Metal1 ;
        RECT 3.655 3.015 3.885 4.360 ;
        RECT 3.655 2.785 4.900 3.015 ;
        RECT 4.670 1.985 4.900 2.785 ;
        RECT 4.670 1.755 6.540 1.985 ;
        RECT 4.670 1.140 4.955 1.755 ;
        RECT 6.310 1.590 6.540 1.755 ;
        RECT 6.310 1.210 7.195 1.590 ;
        RECT 6.965 0.715 7.195 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.840 5.490 ;
        RECT 0.345 3.550 0.575 4.590 ;
        RECT 6.865 3.550 7.095 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 8.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.525 ;
        RECT 2.485 0.450 2.715 1.525 ;
        RECT 0.000 -0.450 7.840 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 1.755 3.175 1.985 ;
        RECT 1.365 0.715 1.595 1.755 ;
        RECT 2.945 0.910 3.175 1.755 ;
        RECT 3.605 0.910 3.835 1.525 ;
        RECT 5.845 0.910 6.075 1.525 ;
        RECT 2.945 0.680 6.075 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai33_1
MACRO gf180mcu_fd_sc_mcu9t5v0__oai33_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai33_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.590 2.280 9.930 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.550 2.050 8.890 2.500 ;
        RECT 10.160 2.270 12.220 2.500 ;
        RECT 10.160 2.050 10.390 2.270 ;
        RECT 8.550 1.820 10.390 2.050 ;
        RECT 8.550 1.770 8.810 1.820 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.430 2.940 13.235 3.170 ;
        RECT 7.430 2.215 7.735 2.940 ;
        RECT 13.005 2.215 13.235 2.940 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.920 2.270 3.260 2.710 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.990 2.270 2.650 2.500 ;
        RECT 2.390 2.000 2.650 2.270 ;
        RECT 3.490 2.270 5.500 2.500 ;
        RECT 3.490 2.000 3.720 2.270 ;
        RECT 2.390 1.770 3.720 2.000 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.940 5.960 3.170 ;
        RECT 0.710 2.215 1.015 2.940 ;
        RECT 5.730 2.500 5.960 2.940 ;
        RECT 5.730 2.270 6.620 2.500 ;
    END
  END B3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.328400 ;
    PORT
      LAYER Metal1 ;
        RECT 3.655 3.630 3.885 4.360 ;
        RECT 10.275 3.630 10.505 4.360 ;
        RECT 3.655 3.400 13.695 3.630 ;
        RECT 13.465 1.590 13.695 3.400 ;
        RECT 10.230 1.480 13.695 1.590 ;
        RECT 8.030 1.250 13.695 1.480 ;
        RECT 10.230 1.140 10.555 1.250 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.560 5.490 ;
        RECT 0.345 3.860 0.575 4.590 ;
        RECT 6.915 3.860 7.145 4.590 ;
        RECT 13.585 3.860 13.815 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.455 ;
        RECT 3.605 0.450 3.835 1.000 ;
        RECT 5.845 0.450 6.075 1.565 ;
        RECT 0.000 -0.450 14.560 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.685 2.160 1.915 ;
        RECT 0.245 0.845 0.475 1.685 ;
        RECT 1.930 1.540 2.160 1.685 ;
        RECT 4.725 1.795 7.195 2.025 ;
        RECT 4.725 1.540 4.955 1.795 ;
        RECT 1.930 1.310 4.955 1.540 ;
        RECT 1.930 0.730 2.715 1.310 ;
        RECT 4.725 0.730 4.955 1.310 ;
        RECT 6.965 1.020 7.195 1.795 ;
        RECT 6.965 0.910 9.435 1.020 ;
        RECT 11.445 0.910 13.915 1.020 ;
        RECT 6.965 0.680 13.915 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai33_2
MACRO gf180mcu_fd_sc_mcu9t5v0__oai33_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai33_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.325 2.190 17.850 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.120 2.495 27.195 2.725 ;
        RECT 19.120 2.270 19.460 2.495 ;
        RECT 21.990 2.270 22.820 2.495 ;
        RECT 26.965 2.215 27.195 2.495 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.690 2.040 20.580 2.265 ;
        RECT 24.720 2.040 25.060 2.265 ;
        RECT 19.690 1.810 25.060 2.040 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.325 2.190 12.795 2.710 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.820 2.650 7.030 2.880 ;
        RECT 0.820 2.190 1.160 2.650 ;
        RECT 4.040 2.270 4.380 2.650 ;
        RECT 6.800 2.500 7.030 2.650 ;
        RECT 6.800 2.270 8.860 2.500 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.000 2.170 2.420 ;
        RECT 4.610 2.190 6.570 2.420 ;
        RECT 4.610 2.000 4.840 2.190 ;
        RECT 1.830 1.770 4.840 2.000 ;
    END
  END B3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 8.382299 ;
    PORT
      LAYER Metal1 ;
        RECT 10.325 3.185 10.555 3.830 ;
        RECT 12.565 3.185 13.850 3.830 ;
        RECT 15.325 3.185 15.555 3.460 ;
        RECT 17.515 3.185 17.745 3.460 ;
        RECT 10.325 2.955 27.655 3.185 ;
        RECT 27.425 1.530 27.655 2.955 ;
        RECT 15.270 1.300 27.655 1.530 ;
        RECT 17.510 1.140 17.850 1.300 ;
        RECT 19.750 1.140 20.090 1.300 ;
        RECT 21.990 1.140 22.330 1.300 ;
        RECT 24.230 1.140 24.570 1.300 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 28.560 5.490 ;
        RECT 2.385 3.580 2.615 4.590 ;
        RECT 6.865 3.580 7.095 4.590 ;
        RECT 20.875 4.150 21.105 4.590 ;
        RECT 25.355 3.875 25.585 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 28.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 28.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.070 ;
        RECT 3.605 0.450 3.835 1.070 ;
        RECT 5.845 0.450 6.075 1.070 ;
        RECT 8.085 0.450 8.315 1.070 ;
        RECT 10.325 0.450 10.555 1.070 ;
        RECT 12.565 0.450 12.795 1.070 ;
        RECT 0.000 -0.450 28.560 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 7.325 4.060 13.870 4.290 ;
        RECT 0.295 3.350 0.525 3.930 ;
        RECT 4.675 3.350 4.905 3.930 ;
        RECT 7.325 3.350 7.555 4.060 ;
        RECT 11.345 3.480 11.575 4.060 ;
        RECT 14.305 3.690 23.345 3.920 ;
        RECT 14.305 3.480 14.535 3.690 ;
        RECT 16.445 3.480 16.675 3.690 ;
        RECT 23.115 3.645 23.345 3.690 ;
        RECT 27.545 3.645 27.775 4.225 ;
        RECT 23.115 3.415 27.775 3.645 ;
        RECT 0.295 3.120 7.555 3.350 ;
        RECT 0.245 1.310 14.430 1.540 ;
        RECT 0.245 0.730 0.475 1.310 ;
        RECT 2.485 0.730 2.715 1.310 ;
        RECT 4.725 0.730 4.955 1.310 ;
        RECT 6.965 0.730 7.195 1.310 ;
        RECT 9.205 0.730 9.435 1.310 ;
        RECT 11.445 0.730 11.675 1.310 ;
        RECT 14.200 1.070 14.430 1.310 ;
        RECT 14.200 0.910 16.675 1.070 ;
        RECT 18.630 0.910 18.970 1.015 ;
        RECT 20.870 0.910 21.210 1.015 ;
        RECT 23.110 0.910 23.450 1.015 ;
        RECT 25.405 0.910 27.875 1.070 ;
        RECT 14.200 0.680 27.875 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai33_4
MACRO gf180mcu_fd_sc_mcu9t5v0__oai211_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai211_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.270 2.170 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.215 1.015 2.710 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 2.270 3.290 2.710 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.990 2.270 4.330 2.710 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.498800 ;
    PORT
      LAYER Metal1 ;
        RECT 2.385 3.320 2.615 4.360 ;
        RECT 4.605 3.320 4.835 4.360 ;
        RECT 1.270 3.090 4.835 3.320 ;
        RECT 1.270 1.140 1.595 3.090 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.600 5.490 ;
        RECT 0.345 3.550 0.575 4.590 ;
        RECT 3.585 3.550 3.815 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 4.605 0.450 4.835 1.655 ;
        RECT 0.000 -0.450 5.600 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 0.910 0.475 1.655 ;
        RECT 2.485 0.910 2.715 1.655 ;
        RECT 0.245 0.680 2.715 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai211_1
MACRO gf180mcu_fd_sc_mcu9t5v0__oai211_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai211_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.795 2.215 2.090 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.200 2.940 2.620 3.170 ;
        RECT 1.200 2.270 1.540 2.940 ;
        RECT 2.390 2.710 2.620 2.940 ;
        RECT 2.390 2.270 4.330 2.710 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.330 2.940 8.535 3.170 ;
        RECT 5.330 2.270 5.670 2.940 ;
        RECT 6.870 2.215 8.535 2.940 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.230 2.270 6.570 2.710 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.025800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.865 4.070 2.665 4.360 ;
        RECT 0.865 3.580 1.095 4.070 ;
        RECT 0.740 3.375 1.095 3.580 ;
        RECT 2.435 3.630 2.665 4.070 ;
        RECT 5.825 3.630 6.055 4.360 ;
        RECT 7.865 3.630 8.095 4.360 ;
        RECT 2.435 3.400 8.095 3.630 ;
        RECT 0.740 1.570 0.970 3.375 ;
        RECT 0.740 1.340 3.890 1.570 ;
        RECT 0.740 1.140 1.595 1.340 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 9.520 5.490 ;
        RECT 0.345 3.860 0.575 4.590 ;
        RECT 4.625 3.860 4.855 4.590 ;
        RECT 6.845 3.860 7.075 4.590 ;
        RECT 8.885 3.860 9.115 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 6.845 0.450 7.075 1.525 ;
        RECT 0.000 -0.450 9.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 4.725 1.755 9.115 1.985 ;
        RECT 0.245 0.910 0.475 1.580 ;
        RECT 4.725 1.110 4.955 1.755 ;
        RECT 2.485 0.910 4.955 1.110 ;
        RECT 0.245 0.680 4.955 0.910 ;
        RECT 8.885 0.770 9.115 1.755 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai211_2
MACRO gf180mcu_fd_sc_mcu9t5v0__oai211_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai211_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.060 2.390 3.770 2.620 ;
        RECT 3.510 2.100 3.770 2.390 ;
        RECT 4.560 2.390 6.620 2.620 ;
        RECT 4.560 2.100 4.790 2.390 ;
        RECT 3.510 1.870 4.790 2.100 ;
        RECT 3.510 1.770 3.770 1.870 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.870 2.850 7.080 3.080 ;
        RECT 0.870 2.390 1.210 2.850 ;
        RECT 4.070 2.330 4.330 2.850 ;
        RECT 6.850 2.620 7.080 2.850 ;
        RECT 6.850 2.390 8.810 2.620 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.670 2.850 15.470 3.080 ;
        RECT 9.670 2.330 9.955 2.850 ;
        RECT 12.875 2.335 13.105 2.850 ;
        RECT 15.240 2.620 15.470 2.850 ;
        RECT 15.240 2.390 17.150 2.620 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.850 2.390 12.500 2.620 ;
        RECT 12.270 2.155 12.500 2.390 ;
        RECT 13.335 2.390 15.010 2.620 ;
        RECT 12.270 2.000 12.730 2.155 ;
        RECT 13.335 2.000 13.565 2.390 ;
        RECT 12.330 1.770 13.565 2.000 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.960100 ;
    PORT
      LAYER Metal1 ;
        RECT 2.485 3.540 2.715 4.360 ;
        RECT 6.915 3.540 7.145 4.360 ;
        RECT 10.305 3.540 10.535 4.120 ;
        RECT 12.345 3.830 12.575 4.360 ;
        RECT 11.910 3.540 12.575 3.830 ;
        RECT 14.385 3.540 14.615 4.345 ;
        RECT 16.425 3.540 16.655 4.360 ;
        RECT 0.410 3.310 16.655 3.540 ;
        RECT 0.410 1.950 0.640 3.310 ;
        RECT 0.410 1.720 3.280 1.950 ;
        RECT 1.365 1.140 1.595 1.720 ;
        RECT 3.050 1.540 3.280 1.720 ;
        RECT 5.980 1.600 8.315 1.830 ;
        RECT 5.980 1.580 6.210 1.600 ;
        RECT 3.990 1.540 6.210 1.580 ;
        RECT 3.050 1.350 6.210 1.540 ;
        RECT 3.050 1.140 4.120 1.350 ;
        RECT 5.845 1.140 6.210 1.350 ;
        RECT 8.085 1.140 8.315 1.600 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.920 5.490 ;
        RECT 0.345 3.770 0.575 4.590 ;
        RECT 4.675 3.770 4.905 4.590 ;
        RECT 9.105 3.770 9.335 4.590 ;
        RECT 11.325 3.770 11.555 4.590 ;
        RECT 13.365 3.770 13.595 4.590 ;
        RECT 15.405 3.770 15.635 4.590 ;
        RECT 17.445 3.770 17.675 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 18.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 11.325 0.450 11.555 1.265 ;
        RECT 15.405 0.450 15.635 1.490 ;
        RECT 0.000 -0.450 17.920 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 9.205 1.540 12.100 1.725 ;
        RECT 13.795 1.720 17.675 1.950 ;
        RECT 13.795 1.540 14.025 1.720 ;
        RECT 9.205 1.495 14.025 1.540 ;
        RECT 0.245 0.910 0.475 1.490 ;
        RECT 2.430 0.910 2.770 0.965 ;
        RECT 4.670 0.910 5.010 0.965 ;
        RECT 6.910 0.910 7.250 0.965 ;
        RECT 9.205 0.910 9.435 1.495 ;
        RECT 11.870 1.310 14.025 1.495 ;
        RECT 0.245 0.680 9.435 0.910 ;
        RECT 13.365 0.680 13.595 1.310 ;
        RECT 17.445 0.680 17.675 1.720 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai211_4
MACRO gf180mcu_fd_sc_mcu9t5v0__oai221_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai221_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.190 1.770 5.455 2.555 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.070 2.215 4.435 2.710 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.150 2.090 2.710 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 1.015 2.555 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 2.270 3.290 2.710 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.661600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.565 3.320 2.795 4.360 ;
        RECT 5.805 3.320 6.035 4.360 ;
        RECT 2.565 3.090 6.035 3.320 ;
        RECT 4.665 1.590 4.895 3.090 ;
        RECT 4.630 1.480 4.895 1.590 ;
        RECT 4.630 1.140 5.015 1.480 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 6.720 5.490 ;
        RECT 0.345 3.550 0.575 4.590 ;
        RECT 3.585 3.550 3.815 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.150 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.150 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.070 ;
        RECT 0.000 -0.450 6.720 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.310 2.715 1.540 ;
        RECT 0.245 0.730 0.475 1.310 ;
        RECT 2.485 0.730 2.715 1.310 ;
        RECT 3.665 0.910 3.895 1.540 ;
        RECT 5.905 0.910 6.135 1.540 ;
        RECT 3.665 0.680 6.135 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai221_1
MACRO gf180mcu_fd_sc_mcu9t5v0__oai221_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai221_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.320 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.530 2.890 9.305 3.270 ;
        RECT 7.530 2.215 7.760 2.890 ;
        RECT 9.075 2.500 9.305 2.890 ;
        RECT 9.075 2.270 11.140 2.500 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.990 2.215 8.845 2.555 ;
        RECT 7.990 1.770 8.250 2.215 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 2.150 3.210 2.710 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.270 2.940 4.805 3.170 ;
        RECT 2.270 2.555 2.500 2.940 ;
        RECT 1.210 2.325 2.500 2.555 ;
        RECT 4.575 2.555 4.805 2.940 ;
        RECT 1.210 1.830 2.165 2.325 ;
        RECT 4.575 2.215 5.425 2.555 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.980 3.580 5.265 3.630 ;
        RECT 0.710 3.400 5.265 3.580 ;
        RECT 0.710 3.350 2.125 3.400 ;
        RECT 0.710 1.770 0.970 3.350 ;
        RECT 5.035 3.015 5.265 3.400 ;
        RECT 5.035 2.785 6.625 3.015 ;
        RECT 6.395 2.215 6.625 2.785 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.216500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.295 4.040 0.525 4.360 ;
        RECT 3.535 4.090 3.765 4.360 ;
        RECT 1.690 4.040 5.725 4.090 ;
        RECT 0.295 3.860 5.725 4.040 ;
        RECT 0.295 3.810 1.835 3.860 ;
        RECT 5.495 3.780 5.725 3.860 ;
        RECT 6.975 3.780 7.205 4.360 ;
        RECT 5.495 3.550 11.665 3.780 ;
        RECT 10.790 2.890 11.665 3.550 ;
        RECT 11.435 1.985 11.665 2.890 ;
        RECT 8.480 1.755 11.665 1.985 ;
        RECT 8.480 1.540 8.710 1.755 ;
        RECT 8.120 1.310 8.710 1.540 ;
        RECT 10.415 1.140 10.645 1.755 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 12.320 5.490 ;
        RECT 1.315 4.270 1.545 4.590 ;
        RECT 5.955 4.020 6.185 4.590 ;
        RECT 9.245 4.020 9.475 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 12.750 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.750 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.460 0.450 2.800 0.640 ;
        RECT 4.700 0.450 5.040 0.640 ;
        RECT 0.000 -0.450 12.320 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.100 0.475 1.525 ;
        RECT 1.340 1.330 6.160 1.560 ;
        RECT 7.055 1.100 7.285 1.190 ;
        RECT 0.245 0.910 7.285 1.100 ;
        RECT 9.295 0.910 9.525 1.525 ;
        RECT 11.535 0.910 11.765 1.525 ;
        RECT 0.245 0.870 11.765 0.910 ;
        RECT 0.245 0.715 0.475 0.870 ;
        RECT 7.055 0.680 11.765 0.870 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai221_2
MACRO gf180mcu_fd_sc_mcu9t5v0__oai221_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai221_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.080 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.030 3.040 21.190 3.270 ;
        RECT 15.030 2.270 15.370 3.040 ;
        RECT 19.140 2.890 21.190 3.040 ;
        RECT 19.140 2.215 19.370 2.890 ;
        RECT 20.960 2.500 21.190 2.890 ;
        RECT 20.960 2.270 22.970 2.500 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 17.270 2.270 17.770 2.500 ;
        RECT 17.510 1.985 17.770 2.270 ;
        RECT 19.600 2.270 20.730 2.500 ;
        RECT 19.600 1.985 19.830 2.270 ;
        RECT 17.510 1.755 19.830 1.985 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.870 2.730 7.080 2.960 ;
        RECT 0.870 2.270 1.210 2.730 ;
        RECT 4.070 2.270 4.410 2.730 ;
        RECT 6.850 2.500 7.080 2.730 ;
        RECT 6.850 2.270 8.860 2.500 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.060 2.270 3.630 2.500 ;
        RECT 3.400 2.175 3.630 2.270 ;
        RECT 4.640 2.270 6.620 2.500 ;
        RECT 3.400 2.040 3.860 2.175 ;
        RECT 4.640 2.040 4.870 2.270 ;
        RECT 3.400 2.020 4.870 2.040 ;
        RECT 3.460 1.770 4.870 2.020 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.990 2.270 13.570 2.710 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 10.615000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.345 3.420 0.575 4.360 ;
        RECT 4.675 3.730 4.905 4.360 ;
        RECT 9.155 3.730 9.385 4.360 ;
        RECT 12.165 3.730 12.395 4.360 ;
        RECT 14.305 3.730 14.535 4.360 ;
        RECT 18.570 3.730 19.065 4.360 ;
        RECT 23.265 3.730 23.495 4.360 ;
        RECT 4.675 3.500 23.495 3.730 ;
        RECT 4.675 3.420 4.905 3.500 ;
        RECT 0.345 3.190 4.905 3.420 ;
        RECT 23.200 1.970 23.495 3.500 ;
        RECT 20.060 1.740 23.495 1.970 ;
        RECT 20.060 1.520 20.290 1.740 ;
        RECT 15.525 1.290 20.290 1.520 ;
        RECT 15.525 1.140 15.755 1.290 ;
        RECT 17.710 1.140 18.050 1.290 ;
        RECT 20.005 1.140 20.290 1.290 ;
        RECT 22.245 1.140 22.475 1.740 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 24.080 5.490 ;
        RECT 2.435 3.650 2.665 4.590 ;
        RECT 6.915 3.960 7.145 4.590 ;
        RECT 10.945 3.960 11.175 4.590 ;
        RECT 13.185 3.960 13.415 4.590 ;
        RECT 16.595 3.960 16.825 4.590 ;
        RECT 21.075 3.960 21.305 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 24.510 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 24.510 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.510 ;
        RECT 2.485 0.450 2.715 1.510 ;
        RECT 4.725 0.450 4.955 1.040 ;
        RECT 6.965 0.450 7.195 1.040 ;
        RECT 9.205 0.450 9.435 1.040 ;
        RECT 0.000 -0.450 24.080 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 1.740 3.175 1.970 ;
        RECT 1.365 0.700 1.595 1.740 ;
        RECT 2.945 1.510 3.175 1.740 ;
        RECT 2.945 1.280 13.515 1.510 ;
        RECT 3.605 0.700 3.835 1.280 ;
        RECT 5.845 0.700 6.075 1.280 ;
        RECT 8.085 0.700 8.315 1.280 ;
        RECT 10.990 1.140 11.330 1.280 ;
        RECT 13.285 1.140 13.515 1.280 ;
        RECT 9.925 0.910 10.155 1.040 ;
        RECT 12.110 0.910 12.450 0.985 ;
        RECT 14.350 0.910 14.690 0.985 ;
        RECT 16.590 0.910 16.930 0.985 ;
        RECT 18.830 0.910 19.170 0.985 ;
        RECT 21.125 0.910 21.355 1.510 ;
        RECT 23.365 0.910 23.595 1.510 ;
        RECT 9.925 0.680 23.595 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai221_4
MACRO gf180mcu_fd_sc_mcu9t5v0__oai222_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai222_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.400 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.870 2.270 7.290 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 2.270 6.180 2.710 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 1.770 3.980 2.500 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.630 2.270 5.050 2.710 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.150 2.090 2.710 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.215 1.015 2.710 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.943800 ;
    PORT
      LAYER Metal1 ;
        RECT 3.255 3.830 3.485 4.360 ;
        RECT 7.585 3.830 7.815 4.360 ;
        RECT 3.255 3.550 7.815 3.830 ;
        RECT 3.255 3.450 6.640 3.550 ;
        RECT 6.410 1.480 6.640 3.450 ;
        RECT 6.410 1.140 6.795 1.480 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 8.400 5.490 ;
        RECT 0.345 3.550 0.575 4.590 ;
        RECT 5.345 4.060 5.575 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 8.830 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.830 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.205 ;
        RECT 0.000 -0.450 8.400 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 1.540 3.305 1.665 ;
        RECT 1.365 1.435 4.555 1.540 ;
        RECT 1.365 0.680 1.595 1.435 ;
        RECT 3.100 1.310 4.555 1.435 ;
        RECT 4.325 1.140 4.555 1.310 ;
        RECT 3.150 0.910 3.490 0.965 ;
        RECT 5.445 0.910 5.675 1.490 ;
        RECT 7.685 0.910 7.915 1.490 ;
        RECT 3.150 0.680 7.915 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai222_1
MACRO gf180mcu_fd_sc_mcu9t5v0__oai222_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai222_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.120 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.605 2.940 12.500 3.170 ;
        RECT 10.605 2.215 10.835 2.940 ;
        RECT 12.270 2.710 12.500 2.940 ;
        RECT 12.270 2.215 14.005 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.350 2.215 11.715 2.710 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.190 3.040 9.525 3.270 ;
        RECT 5.190 2.215 6.165 3.040 ;
        RECT 9.295 2.215 9.525 3.040 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.870 2.215 7.285 2.710 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.925 2.785 4.330 3.015 ;
        RECT 0.925 2.215 1.155 2.785 ;
        RECT 4.070 1.770 4.330 2.785 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.090 2.555 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.570000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.345 3.550 0.575 4.360 ;
        RECT 4.675 3.730 4.905 4.360 ;
        RECT 8.490 4.130 10.105 4.360 ;
        RECT 8.490 3.730 8.870 4.130 ;
        RECT 4.675 3.550 8.870 3.730 ;
        RECT 0.345 3.500 8.870 3.550 ;
        RECT 9.875 3.630 10.105 4.130 ;
        RECT 14.355 3.630 14.585 4.360 ;
        RECT 0.345 3.320 4.900 3.500 ;
        RECT 9.875 3.400 14.585 3.630 ;
        RECT 14.355 1.950 14.585 3.400 ;
        RECT 11.045 1.720 14.585 1.950 ;
        RECT 11.045 1.140 11.275 1.720 ;
        RECT 13.285 1.140 13.515 1.720 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 15.120 5.490 ;
        RECT 2.435 3.780 2.665 4.590 ;
        RECT 7.635 3.960 7.865 4.590 ;
        RECT 12.115 3.860 12.345 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 15.550 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 15.550 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.655 ;
        RECT 2.485 0.450 2.715 0.695 ;
        RECT 4.725 0.450 4.955 0.695 ;
        RECT 0.000 -0.450 15.120 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 1.140 9.035 1.540 ;
        RECT 1.365 0.925 3.835 1.140 ;
        RECT 1.365 0.730 1.595 0.925 ;
        RECT 3.605 0.730 3.835 0.925 ;
        RECT 9.925 0.910 10.155 1.575 ;
        RECT 12.165 0.910 12.395 1.490 ;
        RECT 14.405 0.910 14.635 1.490 ;
        RECT 5.390 0.680 14.635 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai222_2
MACRO gf180mcu_fd_sc_mcu9t5v0__oai222_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai222_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.190 2.000 19.660 2.500 ;
        RECT 22.685 2.000 22.915 2.145 ;
        RECT 27.165 2.000 27.395 2.555 ;
        RECT 19.190 1.770 27.395 2.000 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 21.700 2.480 25.260 2.710 ;
        RECT 21.700 2.270 22.040 2.480 ;
        RECT 23.110 2.270 25.260 2.480 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.605 3.040 18.540 3.270 ;
        RECT 10.605 2.890 14.060 3.040 ;
        RECT 10.605 2.215 10.835 2.890 ;
        RECT 13.720 2.270 14.060 2.890 ;
        RECT 18.200 2.270 18.540 3.040 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.740 2.270 13.290 2.500 ;
        RECT 13.030 2.000 13.290 2.270 ;
        RECT 14.290 2.270 16.250 2.500 ;
        RECT 14.290 2.000 14.520 2.270 ;
        RECT 13.030 1.770 14.520 2.000 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.875 2.785 7.080 3.015 ;
        RECT 0.875 2.215 1.105 2.785 ;
        RECT 4.040 2.270 4.380 2.785 ;
        RECT 6.850 2.500 7.080 2.785 ;
        RECT 6.850 2.270 8.860 2.500 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.165 2.215 3.770 2.555 ;
        RECT 3.510 2.000 3.770 2.215 ;
        RECT 4.610 2.270 6.620 2.500 ;
        RECT 4.610 2.000 4.840 2.270 ;
        RECT 3.510 1.770 4.840 2.000 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 11.529600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.295 3.475 0.525 4.360 ;
        RECT 4.675 3.550 4.905 4.360 ;
        RECT 9.155 3.730 9.385 4.360 ;
        RECT 12.970 3.730 14.585 4.360 ;
        RECT 18.835 3.730 19.065 4.360 ;
        RECT 9.155 3.550 19.065 3.730 ;
        RECT 4.675 3.500 19.065 3.550 ;
        RECT 4.675 3.475 9.380 3.500 ;
        RECT 0.295 3.245 9.380 3.475 ;
        RECT 18.835 3.320 19.065 3.500 ;
        RECT 23.265 3.320 23.495 4.360 ;
        RECT 27.745 3.320 27.975 4.360 ;
        RECT 18.835 3.090 27.975 3.320 ;
        RECT 27.745 1.515 27.975 3.090 ;
        RECT 20.005 1.285 27.975 1.515 ;
        RECT 20.005 1.140 20.235 1.285 ;
        RECT 22.190 1.140 22.530 1.285 ;
        RECT 24.430 1.140 24.770 1.285 ;
        RECT 26.670 1.140 27.010 1.285 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 28.560 5.490 ;
        RECT 2.435 3.705 2.665 4.590 ;
        RECT 6.915 3.780 7.145 4.590 ;
        RECT 12.115 3.960 12.345 4.590 ;
        RECT 16.595 3.960 16.825 4.590 ;
        RECT 21.075 3.550 21.305 4.590 ;
        RECT 25.555 3.550 25.785 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 28.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 28.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.525 ;
        RECT 2.485 0.450 2.715 1.525 ;
        RECT 4.725 0.450 4.955 1.055 ;
        RECT 6.965 0.450 7.195 1.525 ;
        RECT 9.205 0.450 9.435 1.525 ;
        RECT 0.000 -0.450 28.560 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 1.755 3.280 1.985 ;
        RECT 1.365 0.715 1.595 1.755 ;
        RECT 3.050 1.525 3.280 1.755 ;
        RECT 5.845 1.755 11.220 1.985 ;
        RECT 5.845 1.525 6.075 1.755 ;
        RECT 3.050 1.295 6.075 1.525 ;
        RECT 3.605 0.715 3.835 1.295 ;
        RECT 5.845 0.715 6.075 1.295 ;
        RECT 8.085 0.715 8.315 1.755 ;
        RECT 9.925 0.910 10.155 1.525 ;
        RECT 10.990 1.520 11.220 1.755 ;
        RECT 15.580 1.755 17.995 1.985 ;
        RECT 15.580 1.520 15.810 1.755 ;
        RECT 10.990 1.290 15.810 1.520 ;
        RECT 10.990 1.140 11.275 1.290 ;
        RECT 13.230 1.140 13.570 1.290 ;
        RECT 15.525 1.140 15.810 1.290 ;
        RECT 12.110 0.910 12.450 1.000 ;
        RECT 14.350 0.910 14.690 1.000 ;
        RECT 16.645 0.910 16.875 1.525 ;
        RECT 17.765 1.140 17.995 1.755 ;
        RECT 18.885 0.910 19.115 1.525 ;
        RECT 21.070 0.910 21.410 1.000 ;
        RECT 23.310 0.910 23.650 1.000 ;
        RECT 25.550 0.910 25.890 1.000 ;
        RECT 27.845 0.910 28.075 1.055 ;
        RECT 9.925 0.680 28.075 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai222_4
MACRO gf180mcu_fd_sc_mcu9t5v0__or2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.853500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.215 1.070 3.270 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.853500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.210 2.090 2.555 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.800 1.590 4.130 4.360 ;
        RECT 3.510 1.210 4.130 1.590 ;
        RECT 3.900 0.680 4.130 1.210 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 4.480 5.490 ;
        RECT 2.780 3.790 3.010 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 4.910 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 0.450 0.530 0.995 ;
        RECT 2.780 0.450 3.010 0.995 ;
        RECT 0.000 -0.450 4.480 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.845 2.550 4.075 ;
        RECT 2.320 2.500 2.550 3.845 ;
        RECT 2.320 2.270 3.505 2.500 ;
        RECT 2.320 0.940 2.550 2.270 ;
        RECT 1.365 0.710 2.550 0.940 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or2_1
MACRO gf180mcu_fd_sc_mcu9t5v0__or2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.270 1.070 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.795 2.215 2.090 2.710 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.729500 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 0.680 3.835 4.360 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 5.600 5.490 ;
        RECT 2.435 3.550 2.665 4.590 ;
        RECT 4.625 3.550 4.855 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.030 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 0.000 -0.450 5.600 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.320 0.575 4.360 ;
        RECT 0.345 3.090 3.205 3.320 ;
        RECT 2.975 1.950 3.205 3.090 ;
        RECT 1.365 1.720 3.205 1.950 ;
        RECT 1.365 0.680 1.595 1.720 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or2_2
MACRO gf180mcu_fd_sc_mcu9t5v0__or2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 2.270 2.140 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.870 2.940 4.275 3.170 ;
        RECT 0.870 2.270 1.210 2.940 ;
        RECT 2.390 2.215 4.275 2.940 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.550500 ;
    PORT
      LAYER Metal1 ;
        RECT 6.085 3.320 6.315 4.360 ;
        RECT 8.175 3.320 8.405 4.360 ;
        RECT 6.085 3.090 8.405 3.320 ;
        RECT 7.620 1.590 7.850 3.090 ;
        RECT 5.985 1.490 7.850 1.590 ;
        RECT 5.985 1.210 8.455 1.490 ;
        RECT 5.985 0.680 6.215 1.210 ;
        RECT 8.225 0.680 8.455 1.210 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 10.080 5.490 ;
        RECT 0.345 3.550 0.575 4.590 ;
        RECT 4.965 3.550 5.195 4.590 ;
        RECT 7.105 3.550 7.335 4.590 ;
        RECT 9.245 3.550 9.475 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 10.510 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.490 ;
        RECT 2.485 0.450 2.715 1.490 ;
        RECT 4.725 0.450 4.955 1.490 ;
        RECT 7.105 0.450 7.335 0.980 ;
        RECT 9.345 0.450 9.575 1.490 ;
        RECT 0.000 -0.450 10.080 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.535 3.630 2.765 4.360 ;
        RECT 2.535 3.400 4.735 3.630 ;
        RECT 4.505 2.500 4.735 3.400 ;
        RECT 4.505 2.270 7.390 2.500 ;
        RECT 4.505 1.970 4.735 2.270 ;
        RECT 1.365 1.740 4.735 1.970 ;
        RECT 1.365 0.680 1.595 1.740 ;
        RECT 3.605 0.680 3.835 1.740 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or2_4
MACRO gf180mcu_fd_sc_mcu9t5v0__or3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.160 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.772500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.785 2.150 1.015 2.555 ;
        RECT 0.150 1.770 1.015 2.150 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.772500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.090 2.555 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.772500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 2.215 3.335 2.710 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.045 0.680 5.450 4.360 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 6.160 5.490 ;
        RECT 4.025 3.790 4.255 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 6.590 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.590 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 0.860 ;
        RECT 3.785 0.450 4.015 0.860 ;
        RECT 0.000 -0.450 6.160 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.290 3.845 3.795 4.075 ;
        RECT 3.565 2.500 3.795 3.845 ;
        RECT 3.565 2.270 4.750 2.500 ;
        RECT 3.565 1.320 3.795 2.270 ;
        RECT 0.245 1.090 3.795 1.320 ;
        RECT 0.245 0.680 0.475 1.090 ;
        RECT 2.485 0.680 2.715 1.090 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or3_1
MACRO gf180mcu_fd_sc_mcu9t5v0__or3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.545000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.270 1.070 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.545000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.795 2.215 2.090 2.710 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.545000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.915 2.215 3.210 2.710 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.729500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.630 2.890 5.135 4.360 ;
        RECT 4.905 0.680 5.135 2.890 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 6.720 5.490 ;
        RECT 3.555 3.550 3.785 4.590 ;
        RECT 5.925 3.550 6.155 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.150 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.150 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.385 ;
        RECT 3.605 0.450 3.835 1.385 ;
        RECT 6.025 0.450 6.255 1.490 ;
        RECT 0.000 -0.450 6.720 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.320 0.575 4.360 ;
        RECT 0.345 3.090 3.670 3.320 ;
        RECT 3.440 2.555 3.670 3.090 ;
        RECT 3.440 2.215 4.505 2.555 ;
        RECT 3.440 1.845 3.670 2.215 ;
        RECT 0.245 1.615 3.670 1.845 ;
        RECT 0.245 0.680 0.475 1.615 ;
        RECT 2.485 0.680 2.715 1.615 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or3_2
MACRO gf180mcu_fd_sc_mcu9t5v0__or3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.320 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.090000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.920 2.270 3.260 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.090000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.000 2.170 2.500 ;
        RECT 3.490 2.270 5.500 2.500 ;
        RECT 3.490 2.000 3.720 2.270 ;
        RECT 1.830 1.770 3.720 2.000 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.090000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.940 6.570 3.170 ;
        RECT 0.710 2.270 1.070 2.940 ;
        RECT 6.230 2.270 6.570 2.940 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.459000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.315 3.630 8.545 4.360 ;
        RECT 10.455 3.630 10.685 4.360 ;
        RECT 8.315 3.400 10.685 3.630 ;
        RECT 9.900 1.590 10.130 3.400 ;
        RECT 8.265 1.490 10.130 1.590 ;
        RECT 8.265 1.210 10.735 1.490 ;
        RECT 8.265 0.680 8.495 1.210 ;
        RECT 10.505 0.680 10.735 1.210 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 12.320 5.490 ;
        RECT 0.345 3.860 0.575 4.590 ;
        RECT 6.865 3.860 7.095 4.590 ;
        RECT 9.335 3.860 9.565 4.590 ;
        RECT 11.525 3.860 11.755 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 12.750 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.750 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.385 ;
        RECT 2.485 0.450 2.715 0.915 ;
        RECT 4.725 0.450 4.955 0.915 ;
        RECT 6.965 0.450 7.195 0.915 ;
        RECT 9.385 0.450 9.615 0.915 ;
        RECT 11.625 0.450 11.855 1.385 ;
        RECT 0.000 -0.450 12.320 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.655 3.630 3.885 4.360 ;
        RECT 3.655 3.400 7.030 3.630 ;
        RECT 6.800 2.500 7.030 3.400 ;
        RECT 6.800 2.270 9.670 2.500 ;
        RECT 6.800 1.375 7.030 2.270 ;
        RECT 1.365 1.145 7.030 1.375 ;
        RECT 1.365 0.680 1.595 1.145 ;
        RECT 3.605 0.680 3.835 1.145 ;
        RECT 5.845 0.680 6.075 1.145 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or3_4
MACRO gf180mcu_fd_sc_mcu9t5v0__or4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.694500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.785 2.150 1.015 2.555 ;
        RECT 0.150 1.770 1.015 2.150 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.694500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.215 2.555 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.694500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 1.770 3.385 2.555 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.694500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.345 1.590 4.575 2.555 ;
        RECT 4.070 1.210 4.575 1.590 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.285 0.680 6.615 4.360 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.280 5.490 ;
        RECT 5.265 3.790 5.495 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.710 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.015 ;
        RECT 2.665 0.450 2.895 1.015 ;
        RECT 5.265 0.450 5.495 0.940 ;
        RECT 0.000 -0.450 7.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.290 3.845 5.035 4.075 ;
        RECT 4.805 2.500 5.035 3.845 ;
        RECT 4.805 2.270 5.990 2.500 ;
        RECT 1.545 1.245 3.840 1.475 ;
        RECT 1.545 0.680 1.775 1.245 ;
        RECT 3.610 0.930 3.840 1.245 ;
        RECT 4.805 0.930 5.035 2.270 ;
        RECT 3.610 0.700 5.035 0.930 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or4_1
MACRO gf180mcu_fd_sc_mcu9t5v0__or4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.270 1.070 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.090 2.555 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.390 2.270 3.260 2.710 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 2.270 4.380 2.710 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.729500 ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 2.890 6.255 4.360 ;
        RECT 6.025 0.680 6.255 2.890 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 7.840 5.490 ;
        RECT 4.675 3.550 4.905 4.590 ;
        RECT 7.045 3.550 7.275 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 8.270 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.020 ;
        RECT 2.485 0.450 2.715 1.020 ;
        RECT 4.725 0.450 4.955 1.020 ;
        RECT 7.145 0.450 7.375 1.490 ;
        RECT 0.000 -0.450 7.840 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.320 0.575 4.360 ;
        RECT 0.345 3.090 4.840 3.320 ;
        RECT 4.610 2.555 4.840 3.090 ;
        RECT 4.610 2.215 5.625 2.555 ;
        RECT 4.610 1.480 4.840 2.215 ;
        RECT 1.365 1.250 4.840 1.480 ;
        RECT 1.365 0.680 1.595 1.250 ;
        RECT 3.605 0.680 3.835 1.250 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or4_2
MACRO gf180mcu_fd_sc_mcu9t5v0__or4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.035 2.215 4.330 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.440 2.940 4.860 3.170 ;
        RECT 3.440 2.500 3.670 2.940 ;
        RECT 3.060 2.270 3.670 2.500 ;
        RECT 4.630 2.710 4.860 2.940 ;
        RECT 4.630 2.215 6.565 2.710 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.940 1.985 2.280 2.500 ;
        RECT 6.870 2.270 7.740 2.500 ;
        RECT 6.870 1.985 7.130 2.270 ;
        RECT 1.940 1.755 7.130 1.985 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.870 3.400 8.200 3.630 ;
        RECT 0.870 2.890 3.210 3.400 ;
        RECT 0.870 2.270 1.210 2.890 ;
        RECT 7.970 2.500 8.200 3.400 ;
        RECT 7.970 2.270 8.860 2.500 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.550500 ;
    PORT
      LAYER Metal1 ;
        RECT 10.170 3.525 10.735 4.360 ;
        RECT 12.645 3.525 12.875 4.360 ;
        RECT 10.170 3.295 12.875 3.525 ;
        RECT 11.280 1.950 11.835 3.295 ;
        RECT 10.505 1.720 12.975 1.950 ;
        RECT 10.505 0.680 10.735 1.720 ;
        RECT 12.745 0.680 12.975 1.720 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 14.560 5.490 ;
        RECT 0.345 3.755 0.575 4.590 ;
        RECT 9.460 4.275 9.690 4.590 ;
        RECT 11.575 3.755 11.805 4.590 ;
        RECT 13.765 3.755 13.995 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 14.990 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.020 ;
        RECT 2.485 0.450 2.715 1.020 ;
        RECT 4.725 0.450 4.955 1.020 ;
        RECT 6.965 0.450 7.195 1.020 ;
        RECT 9.205 0.450 9.435 1.020 ;
        RECT 11.625 0.450 11.855 1.490 ;
        RECT 13.865 0.450 14.095 1.490 ;
        RECT 0.000 -0.450 14.560 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 4.720 3.860 9.320 4.090 ;
        RECT 9.090 2.500 9.320 3.860 ;
        RECT 9.090 2.270 11.050 2.500 ;
        RECT 9.090 1.480 9.320 2.270 ;
        RECT 1.365 1.250 9.320 1.480 ;
        RECT 1.365 0.680 1.595 1.250 ;
        RECT 3.605 0.680 3.835 1.250 ;
        RECT 5.845 0.680 6.075 1.250 ;
        RECT 8.085 0.680 8.315 1.250 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or4_4
MACRO gf180mcu_fd_sc_mcu9t5v0__sdffq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.630 1.210 4.890 2.520 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.696000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.180 0.915 2.710 ;
        RECT 0.150 1.770 0.410 2.180 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 2.180 2.020 2.710 ;
        RECT 1.270 1.770 1.530 2.180 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.310 1.770 6.835 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.495 2.710 19.725 3.690 ;
        RECT 19.190 1.210 19.725 2.710 ;
        RECT 19.445 0.790 19.725 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 21.280 5.490 ;
        RECT 1.315 3.440 1.545 4.590 ;
        RECT 5.030 3.965 5.370 4.590 ;
        RECT 7.180 3.995 7.520 4.590 ;
        RECT 12.595 3.440 12.825 4.590 ;
        RECT 17.025 3.595 17.255 4.590 ;
        RECT 20.515 3.880 20.745 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.310 21.710 5.470 ;
        RECT -0.430 2.265 0.430 2.310 ;
        RECT 19.210 2.270 21.710 2.310 ;
        RECT 20.850 2.265 21.710 2.270 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 9.270 2.265 17.710 2.310 ;
        RECT -0.430 -0.430 21.710 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.075 ;
        RECT 5.450 0.450 5.790 0.510 ;
        RECT 7.450 0.450 7.790 0.510 ;
        RECT 12.810 0.450 13.150 0.505 ;
        RECT 17.385 0.450 17.615 0.720 ;
        RECT 20.565 0.450 20.795 1.600 ;
        RECT 0.000 -0.450 21.280 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.295 3.210 0.525 4.250 ;
        RECT 3.125 3.735 3.355 4.250 ;
        RECT 9.615 3.735 9.845 3.845 ;
        RECT 3.125 3.505 9.845 3.735 ;
        RECT 3.125 3.440 3.355 3.505 ;
        RECT 0.295 2.980 2.775 3.210 ;
        RECT 2.545 1.535 2.775 2.980 ;
        RECT 6.030 3.045 8.355 3.275 ;
        RECT 6.030 2.935 6.260 3.045 ;
        RECT 8.125 1.540 8.355 3.045 ;
        RECT 0.245 1.305 2.775 1.535 ;
        RECT 0.245 0.790 0.475 1.305 ;
        RECT 6.165 1.200 8.355 1.540 ;
        RECT 8.705 2.520 8.935 3.260 ;
        RECT 8.705 2.180 10.285 2.520 ;
        RECT 8.705 1.220 9.075 2.180 ;
        RECT 10.685 1.950 10.915 4.250 ;
        RECT 14.015 2.980 14.375 4.250 ;
        RECT 12.205 2.750 14.375 2.980 ;
        RECT 12.205 2.180 12.435 2.750 ;
        RECT 13.435 1.950 13.665 2.520 ;
        RECT 10.685 1.720 13.665 1.950 ;
        RECT 3.325 0.970 3.555 1.130 ;
        RECT 9.565 0.970 9.795 1.480 ;
        RECT 10.685 1.360 10.915 1.720 ;
        RECT 14.145 1.360 14.375 2.750 ;
        RECT 15.265 3.365 15.495 4.250 ;
        RECT 15.265 3.135 17.930 3.365 ;
        RECT 15.265 1.360 15.495 3.135 ;
        RECT 15.725 1.020 16.065 2.905 ;
        RECT 16.630 1.545 16.970 2.465 ;
        RECT 17.590 2.235 17.930 3.135 ;
        RECT 18.225 2.520 18.455 4.250 ;
        RECT 18.225 2.290 18.955 2.520 ;
        RECT 18.725 1.545 18.955 2.290 ;
        RECT 16.630 1.315 18.955 1.545 ;
        RECT 3.325 0.740 9.795 0.970 ;
        RECT 11.365 0.735 16.065 1.020 ;
        RECT 11.365 0.680 11.595 0.735 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffq_1
MACRO gf180mcu_fd_sc_mcu9t5v0__sdffq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.400 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.070 2.225 4.835 2.710 ;
        RECT 4.070 1.770 4.330 2.225 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.696000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.225 1.015 2.710 ;
        RECT 0.150 1.770 0.410 2.225 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.135 2.710 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.430 1.770 7.690 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.702050 ;
    PORT
      LAYER Metal1 ;
        RECT 20.790 0.845 21.130 4.250 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 22.400 5.490 ;
        RECT 1.365 3.440 1.595 4.590 ;
        RECT 5.235 3.905 5.465 4.590 ;
        RECT 7.830 3.905 8.170 4.590 ;
        RECT 13.235 3.440 13.465 4.590 ;
        RECT 17.645 3.600 17.875 4.590 ;
        RECT 19.735 3.880 19.965 4.590 ;
        RECT 21.810 3.880 22.040 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 22.830 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 22.830 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.075 ;
        RECT 5.505 0.450 5.735 0.620 ;
        RECT 7.565 0.450 7.795 0.620 ;
        RECT 12.870 0.450 13.100 0.620 ;
        RECT 17.745 0.450 17.975 1.590 ;
        RECT 19.685 0.450 19.915 1.600 ;
        RECT 21.925 0.450 22.155 1.165 ;
        RECT 0.000 -0.450 22.400 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.210 0.575 4.250 ;
        RECT 3.375 4.020 5.005 4.250 ;
        RECT 3.375 3.440 3.605 4.020 ;
        RECT 4.775 3.675 5.005 4.020 ;
        RECT 10.455 3.675 10.685 3.785 ;
        RECT 4.775 3.445 10.685 3.675 ;
        RECT 0.345 2.980 2.895 3.210 ;
        RECT 2.665 1.540 2.895 2.980 ;
        RECT 6.865 2.985 8.555 3.215 ;
        RECT 6.865 2.875 7.095 2.985 ;
        RECT 0.245 1.310 2.895 1.540 ;
        RECT 6.225 1.540 6.455 1.650 ;
        RECT 8.325 1.540 8.555 2.985 ;
        RECT 6.225 1.310 8.555 1.540 ;
        RECT 8.905 2.565 9.135 3.215 ;
        RECT 8.905 2.225 11.125 2.565 ;
        RECT 8.905 1.310 9.135 2.225 ;
        RECT 11.475 1.995 11.705 4.250 ;
        RECT 14.255 3.025 14.485 4.250 ;
        RECT 12.795 2.795 14.485 3.025 ;
        RECT 12.795 2.225 13.025 2.795 ;
        RECT 13.525 1.995 13.755 2.565 ;
        RECT 11.475 1.765 13.755 1.995 ;
        RECT 11.475 1.650 11.705 1.765 ;
        RECT 0.245 0.790 0.475 1.310 ;
        RECT 3.325 1.080 3.555 1.130 ;
        RECT 9.625 1.080 9.855 1.430 ;
        RECT 10.745 1.310 11.705 1.650 ;
        RECT 14.205 1.310 14.485 2.795 ;
        RECT 15.325 3.370 15.555 4.250 ;
        RECT 15.325 3.140 17.895 3.370 ;
        RECT 15.325 1.310 15.555 3.140 ;
        RECT 15.785 1.080 16.015 2.910 ;
        RECT 17.205 2.050 17.435 2.565 ;
        RECT 17.665 2.510 17.895 3.140 ;
        RECT 18.665 2.565 18.895 4.250 ;
        RECT 17.665 2.280 18.370 2.510 ;
        RECT 18.665 2.225 19.410 2.565 ;
        RECT 18.665 2.050 19.095 2.225 ;
        RECT 17.205 1.820 19.095 2.050 ;
        RECT 3.325 0.850 9.855 1.080 ;
        RECT 11.370 0.850 16.015 1.080 ;
        RECT 3.325 0.790 3.555 0.850 ;
        RECT 11.370 0.685 11.710 0.850 ;
        RECT 14.730 0.685 16.015 0.850 ;
        RECT 18.865 0.790 19.095 1.820 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffq_2
MACRO gf180mcu_fd_sc_mcu9t5v0__sdffq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.640 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.070 2.370 4.330 2.710 ;
        RECT 4.070 2.030 4.835 2.370 ;
        RECT 4.070 1.770 4.330 2.030 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.696000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 1.770 0.415 2.710 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.370 0.970 2.710 ;
        RECT 0.710 2.030 2.035 2.370 ;
        RECT 0.710 1.770 0.970 2.030 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.190 1.770 5.625 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.468150 ;
    PORT
      LAYER Metal1 ;
        RECT 20.705 3.645 20.985 4.250 ;
        RECT 22.805 3.645 23.035 4.250 ;
        RECT 20.705 3.415 23.035 3.645 ;
        RECT 20.705 2.150 20.935 3.415 ;
        RECT 20.705 1.920 22.810 2.150 ;
        RECT 20.705 0.845 20.935 1.920 ;
        RECT 22.550 1.655 22.810 1.920 ;
        RECT 22.550 1.210 23.175 1.655 ;
        RECT 22.945 0.845 23.175 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 24.640 5.490 ;
        RECT 1.645 3.440 1.875 4.590 ;
        RECT 5.235 4.135 5.465 4.590 ;
        RECT 5.235 3.905 8.170 4.135 ;
        RECT 13.085 3.440 13.315 4.590 ;
        RECT 17.645 3.550 17.875 4.590 ;
        RECT 19.735 3.875 19.965 4.590 ;
        RECT 21.775 3.875 22.005 4.590 ;
        RECT 23.930 3.875 24.160 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 25.070 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 25.070 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.075 ;
        RECT 5.505 0.450 5.735 0.625 ;
        RECT 7.565 0.450 7.795 0.625 ;
        RECT 12.920 0.450 13.150 0.625 ;
        RECT 17.745 0.450 17.975 1.395 ;
        RECT 19.585 0.450 19.815 1.600 ;
        RECT 21.825 0.450 22.055 1.165 ;
        RECT 24.065 0.450 24.295 1.165 ;
        RECT 0.000 -0.450 24.640 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.625 3.210 0.855 4.250 ;
        RECT 3.405 3.675 3.635 4.250 ;
        RECT 10.290 3.675 10.520 3.785 ;
        RECT 3.405 3.445 10.520 3.675 ;
        RECT 3.405 3.440 3.635 3.445 ;
        RECT 0.625 2.980 3.055 3.210 ;
        RECT 2.825 1.535 3.055 2.980 ;
        RECT 6.865 2.875 8.455 3.215 ;
        RECT 8.225 1.655 8.455 2.875 ;
        RECT 0.245 1.305 3.055 1.535 ;
        RECT 6.225 1.315 8.455 1.655 ;
        RECT 8.905 2.370 9.135 3.215 ;
        RECT 8.905 2.030 11.095 2.370 ;
        RECT 8.905 1.315 9.135 2.030 ;
        RECT 11.325 1.800 11.555 4.250 ;
        RECT 14.205 2.830 14.435 4.250 ;
        RECT 12.645 2.600 14.435 2.830 ;
        RECT 12.645 2.030 12.875 2.600 ;
        RECT 13.525 1.800 13.755 2.370 ;
        RECT 11.325 1.655 13.755 1.800 ;
        RECT 10.745 1.570 13.755 1.655 ;
        RECT 0.245 0.790 0.475 1.305 ;
        RECT 3.325 1.085 3.555 1.130 ;
        RECT 9.625 1.085 9.855 1.435 ;
        RECT 10.745 1.315 11.540 1.570 ;
        RECT 14.205 1.315 14.435 2.600 ;
        RECT 15.325 3.320 15.555 4.250 ;
        RECT 15.325 3.090 17.895 3.320 ;
        RECT 15.325 1.315 15.555 3.090 ;
        RECT 15.785 1.085 16.125 2.860 ;
        RECT 17.205 1.855 17.435 2.370 ;
        RECT 17.665 2.315 17.895 3.090 ;
        RECT 18.735 2.370 18.965 4.250 ;
        RECT 17.665 2.085 18.440 2.315 ;
        RECT 18.735 2.030 20.255 2.370 ;
        RECT 18.735 1.855 19.095 2.030 ;
        RECT 17.205 1.625 19.095 1.855 ;
        RECT 3.325 0.855 9.855 1.085 ;
        RECT 11.370 0.855 16.125 1.085 ;
        RECT 3.325 0.790 3.555 0.855 ;
        RECT 11.370 0.690 11.710 0.855 ;
        RECT 14.730 0.690 16.125 0.855 ;
        RECT 18.865 0.790 19.095 1.625 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffq_4
MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.960 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 2.330 4.330 2.710 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.696000 ;
    PORT
      LAYER Metal1 ;
        RECT 18.630 1.770 18.890 2.710 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.696000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.330 0.970 2.710 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 2.330 2.090 2.710 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.310 2.330 7.130 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 20.870 0.845 21.330 4.250 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 22.960 5.490 ;
        RECT 1.315 3.440 1.545 4.590 ;
        RECT 5.085 3.440 5.315 4.590 ;
        RECT 7.180 4.030 7.520 4.590 ;
        RECT 12.155 3.910 12.385 4.590 ;
        RECT 13.955 3.440 14.185 4.590 ;
        RECT 18.200 3.910 18.430 4.590 ;
        RECT 20.240 3.440 20.470 4.590 ;
        RECT 22.120 3.440 22.350 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 23.390 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 23.390 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.285 ;
        RECT 5.450 0.450 5.680 0.530 ;
        RECT 7.285 0.450 7.515 1.180 ;
        RECT 13.265 0.450 13.495 1.440 ;
        RECT 18.200 0.450 18.430 1.275 ;
        RECT 22.170 0.450 22.400 1.655 ;
        RECT 0.000 -0.450 22.960 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.295 3.210 0.525 4.250 ;
        RECT 3.325 3.210 3.555 4.250 ;
        RECT 5.545 3.525 9.380 3.755 ;
        RECT 5.545 3.210 5.775 3.525 ;
        RECT 0.295 2.980 2.775 3.210 ;
        RECT 3.325 2.980 5.775 3.210 ;
        RECT 6.160 3.010 7.955 3.240 ;
        RECT 2.545 2.100 2.775 2.980 ;
        RECT 4.605 2.100 4.835 2.635 ;
        RECT 7.725 2.100 7.955 3.010 ;
        RECT 8.305 2.580 8.535 3.295 ;
        RECT 10.115 3.095 10.345 4.250 ;
        RECT 11.135 3.670 11.365 4.250 ;
        RECT 13.175 3.670 13.405 4.250 ;
        RECT 11.135 3.440 13.405 3.670 ;
        RECT 10.115 2.865 14.310 3.095 ;
        RECT 8.305 2.390 9.820 2.580 ;
        RECT 0.245 1.870 4.835 2.100 ;
        RECT 6.165 1.870 7.955 2.100 ;
        RECT 8.405 2.350 9.820 2.390 ;
        RECT 0.245 0.945 0.475 1.870 ;
        RECT 3.325 0.990 3.555 1.285 ;
        RECT 6.165 1.210 6.395 1.870 ;
        RECT 6.625 1.410 8.175 1.640 ;
        RECT 3.325 0.980 6.095 0.990 ;
        RECT 6.625 0.980 6.855 1.410 ;
        RECT 3.325 0.760 6.855 0.980 ;
        RECT 6.025 0.750 6.855 0.760 ;
        RECT 7.945 0.910 8.175 1.410 ;
        RECT 8.405 1.140 8.635 2.350 ;
        RECT 9.125 0.910 9.355 1.275 ;
        RECT 10.115 0.945 10.475 2.865 ;
        RECT 10.825 1.900 11.055 2.635 ;
        RECT 11.765 2.360 11.995 2.635 ;
        RECT 13.970 2.590 14.310 2.865 ;
        RECT 14.975 2.435 15.205 4.250 ;
        RECT 14.665 2.360 15.205 2.435 ;
        RECT 11.765 2.205 15.205 2.360 ;
        RECT 15.995 4.020 17.970 4.250 ;
        RECT 11.765 2.130 14.835 2.205 ;
        RECT 10.825 1.670 14.375 1.900 ;
        RECT 7.945 0.680 9.355 0.910 ;
        RECT 14.145 0.925 14.375 1.670 ;
        RECT 14.605 1.155 14.835 2.130 ;
        RECT 15.065 0.925 15.295 1.955 ;
        RECT 15.995 1.440 16.225 4.020 ;
        RECT 15.670 1.210 16.225 1.440 ;
        RECT 16.600 0.925 16.830 3.150 ;
        RECT 17.080 1.155 17.410 3.780 ;
        RECT 17.740 3.680 17.970 4.020 ;
        RECT 18.660 4.010 19.910 4.240 ;
        RECT 18.660 3.680 18.890 4.010 ;
        RECT 17.740 3.450 18.890 3.680 ;
        RECT 19.220 3.170 19.450 3.780 ;
        RECT 17.760 2.940 19.450 3.170 ;
        RECT 17.760 2.295 17.990 2.940 ;
        RECT 19.220 2.065 19.450 2.940 ;
        RECT 19.680 2.295 19.910 4.010 ;
        RECT 20.400 2.065 20.630 2.635 ;
        RECT 19.220 1.835 20.630 2.065 ;
        RECT 20.240 0.945 20.630 1.835 ;
        RECT 14.145 0.695 16.830 0.925 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1
MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 2.330 3.995 3.270 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.144000 ;
    PORT
      LAYER Metal1 ;
        RECT 18.070 2.890 18.890 3.270 ;
        RECT 18.610 1.770 18.890 2.890 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.330 1.530 2.735 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.770 1.830 2.150 2.750 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.310 2.330 7.130 2.735 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.674600 ;
    PORT
      LAYER Metal1 ;
        RECT 21.895 0.840 22.250 4.250 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 23.520 5.490 ;
        RECT 1.365 3.440 1.595 4.590 ;
        RECT 5.085 3.440 5.315 4.590 ;
        RECT 7.175 3.940 7.515 4.590 ;
        RECT 12.030 3.440 12.260 4.590 ;
        RECT 13.770 3.440 14.000 4.590 ;
        RECT 18.070 4.480 18.300 4.590 ;
        RECT 20.330 3.440 20.560 4.590 ;
        RECT 22.915 3.440 23.145 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 23.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 23.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.140 ;
        RECT 5.505 0.450 5.735 0.605 ;
        RECT 7.330 0.450 7.560 1.180 ;
        RECT 13.130 0.450 13.360 1.325 ;
        RECT 17.850 0.450 18.080 1.325 ;
        RECT 20.805 0.450 21.035 1.160 ;
        RECT 23.045 0.450 23.275 1.160 ;
        RECT 0.000 -0.450 23.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.210 0.575 4.250 ;
        RECT 3.125 4.020 4.855 4.250 ;
        RECT 3.125 3.440 3.355 4.020 ;
        RECT 4.625 3.210 4.855 4.020 ;
        RECT 8.970 3.710 9.200 4.250 ;
        RECT 5.545 3.480 9.200 3.710 ;
        RECT 5.545 3.210 5.775 3.480 ;
        RECT 8.970 3.440 9.200 3.480 ;
        RECT 0.345 2.980 2.775 3.210 ;
        RECT 4.625 2.980 5.775 3.210 ;
        RECT 2.545 1.600 2.775 2.980 ;
        RECT 6.155 2.965 7.590 3.195 ;
        RECT 7.360 2.735 7.590 2.965 ;
        RECT 8.250 2.735 8.535 3.250 ;
        RECT 9.990 2.915 10.220 4.250 ;
        RECT 11.010 3.210 11.240 4.250 ;
        RECT 13.050 3.210 13.280 4.250 ;
        RECT 14.790 3.250 15.020 4.250 ;
        RECT 11.010 2.980 13.280 3.210 ;
        RECT 14.250 3.020 15.020 3.250 ;
        RECT 15.810 4.020 20.000 4.250 ;
        RECT 9.990 2.735 10.535 2.915 ;
        RECT 4.650 1.600 4.990 2.735 ;
        RECT 7.360 2.505 7.955 2.735 ;
        RECT 8.250 2.520 9.695 2.735 ;
        RECT 9.990 2.685 13.955 2.735 ;
        RECT 8.450 2.505 9.695 2.520 ;
        RECT 10.310 2.505 13.955 2.685 ;
        RECT 7.360 2.100 7.590 2.505 ;
        RECT 0.245 1.370 4.990 1.600 ;
        RECT 6.210 1.870 7.590 2.100 ;
        RECT 0.245 0.800 0.475 1.370 ;
        RECT 6.210 1.270 6.440 1.870 ;
        RECT 6.670 1.410 8.220 1.640 ;
        RECT 3.270 1.065 3.610 1.085 ;
        RECT 3.270 1.040 6.105 1.065 ;
        RECT 6.670 1.040 6.900 1.410 ;
        RECT 3.270 0.835 6.900 1.040 ;
        RECT 6.000 0.810 6.900 0.835 ;
        RECT 7.990 0.985 8.220 1.410 ;
        RECT 8.450 1.215 8.680 2.505 ;
        RECT 9.190 0.985 9.420 1.325 ;
        RECT 10.310 0.985 10.540 2.505 ;
        RECT 14.250 2.275 14.480 3.020 ;
        RECT 11.535 2.045 14.480 2.275 ;
        RECT 10.835 1.815 11.175 1.960 ;
        RECT 10.835 1.585 14.020 1.815 ;
        RECT 13.790 0.985 14.020 1.585 ;
        RECT 14.250 1.215 14.480 2.045 ;
        RECT 14.790 0.985 15.020 2.790 ;
        RECT 15.810 1.555 16.040 4.020 ;
        RECT 15.390 1.215 16.040 1.555 ;
        RECT 16.270 0.985 16.500 2.790 ;
        RECT 16.730 1.215 17.060 3.780 ;
        RECT 17.410 3.550 19.540 3.780 ;
        RECT 17.410 2.450 17.640 3.550 ;
        RECT 19.310 2.215 19.540 3.550 ;
        RECT 19.770 2.525 20.000 4.020 ;
        RECT 19.310 1.985 20.585 2.215 ;
        RECT 7.990 0.755 9.420 0.985 ;
        RECT 13.790 0.755 16.500 0.985 ;
        RECT 19.990 0.800 20.220 1.985 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2
MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.320 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 2.330 4.490 2.735 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.144000 ;
    PORT
      LAYER Metal1 ;
        RECT 18.630 1.770 18.890 2.790 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 1.175 2.735 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.530 2.735 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.870 1.770 7.400 2.735 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642000 ;
    PORT
      LAYER Metal1 ;
        RECT 22.425 1.620 22.655 4.250 ;
        RECT 24.230 1.620 24.895 4.250 ;
        RECT 22.425 1.390 24.895 1.620 ;
        RECT 22.425 0.840 22.655 1.390 ;
        RECT 24.230 1.210 24.895 1.390 ;
        RECT 24.665 0.840 24.895 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 26.320 5.490 ;
        RECT 1.510 3.440 1.740 4.590 ;
        RECT 5.525 3.440 5.755 4.590 ;
        RECT 7.640 3.940 7.980 4.590 ;
        RECT 12.825 3.450 13.055 4.590 ;
        RECT 14.585 3.440 14.815 4.590 ;
        RECT 18.885 4.350 19.115 4.590 ;
        RECT 20.925 3.440 21.155 4.590 ;
        RECT 23.495 3.440 23.725 4.590 ;
        RECT 25.645 3.440 25.875 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 26.750 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 26.750 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.585 0.450 1.815 1.080 ;
        RECT 5.945 0.450 6.175 0.645 ;
        RECT 7.965 0.450 8.195 0.620 ;
        RECT 13.945 0.450 14.175 1.380 ;
        RECT 18.445 0.450 18.675 1.380 ;
        RECT 21.305 0.450 21.535 1.160 ;
        RECT 23.545 0.450 23.775 1.160 ;
        RECT 25.785 0.450 26.015 1.160 ;
        RECT 0.000 -0.450 26.320 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.490 3.195 0.720 4.250 ;
        RECT 3.765 3.210 3.995 4.250 ;
        RECT 9.765 3.710 9.995 4.250 ;
        RECT 5.985 3.480 9.995 3.710 ;
        RECT 5.985 3.210 6.215 3.480 ;
        RECT 9.765 3.440 9.995 3.480 ;
        RECT 0.490 2.965 3.215 3.195 ;
        RECT 3.765 2.980 6.215 3.210 ;
        RECT 6.620 2.965 7.860 3.195 ;
        RECT 2.985 2.100 3.215 2.965 ;
        RECT 5.145 2.100 5.375 2.750 ;
        RECT 7.630 2.735 7.860 2.965 ;
        RECT 8.715 2.735 8.945 3.250 ;
        RECT 10.785 2.940 11.015 4.250 ;
        RECT 11.805 3.220 12.035 4.250 ;
        RECT 13.845 3.220 14.075 4.250 ;
        RECT 15.605 3.250 15.835 4.250 ;
        RECT 11.805 2.990 14.075 3.220 ;
        RECT 15.065 3.020 15.835 3.250 ;
        RECT 16.625 4.245 18.450 4.250 ;
        RECT 16.625 4.120 18.680 4.245 ;
        RECT 19.245 4.120 20.595 4.160 ;
        RECT 16.625 4.020 20.595 4.120 ;
        RECT 16.625 3.115 16.855 4.020 ;
        RECT 18.400 3.930 20.595 4.020 ;
        RECT 18.400 3.890 19.375 3.930 ;
        RECT 10.785 2.760 11.370 2.940 ;
        RECT 7.630 2.505 8.420 2.735 ;
        RECT 8.715 2.505 10.490 2.735 ;
        RECT 10.785 2.710 14.770 2.760 ;
        RECT 11.145 2.530 14.770 2.710 ;
        RECT 2.985 1.870 5.375 2.100 ;
        RECT 2.985 1.540 3.215 1.870 ;
        RECT 8.190 1.540 8.420 2.505 ;
        RECT 0.245 1.310 3.215 1.540 ;
        RECT 0.245 1.005 0.475 1.310 ;
        RECT 3.765 1.105 3.995 1.345 ;
        RECT 6.570 1.310 8.420 1.540 ;
        RECT 9.305 1.195 9.535 2.505 ;
        RECT 3.765 1.080 6.465 1.105 ;
        RECT 3.765 0.965 9.080 1.080 ;
        RECT 10.025 0.965 10.255 1.380 ;
        RECT 11.145 1.070 11.375 2.530 ;
        RECT 15.065 2.300 15.295 3.020 ;
        RECT 16.185 2.885 16.855 3.115 ;
        RECT 17.525 3.440 17.875 3.780 ;
        RECT 12.370 2.070 15.295 2.300 ;
        RECT 11.670 1.840 12.010 2.015 ;
        RECT 11.670 1.610 14.835 1.840 ;
        RECT 3.765 0.875 10.255 0.965 ;
        RECT 6.360 0.850 10.255 0.875 ;
        RECT 8.855 0.735 10.255 0.850 ;
        RECT 14.605 1.040 14.835 1.610 ;
        RECT 15.065 1.270 15.295 2.070 ;
        RECT 15.605 1.040 15.835 2.790 ;
        RECT 16.185 1.270 16.415 2.885 ;
        RECT 17.065 2.070 17.295 2.790 ;
        RECT 16.865 1.840 17.295 2.070 ;
        RECT 16.865 1.040 17.095 1.840 ;
        RECT 17.525 1.610 17.755 3.440 ;
        RECT 19.905 3.250 20.135 3.700 ;
        RECT 18.005 3.155 20.135 3.250 ;
        RECT 18.005 3.020 20.115 3.155 ;
        RECT 18.005 2.450 18.235 3.020 ;
        RECT 19.885 2.215 20.115 3.020 ;
        RECT 20.365 2.855 20.595 3.930 ;
        RECT 20.345 2.515 20.595 2.855 ;
        RECT 19.885 1.985 21.085 2.215 ;
        RECT 17.325 1.270 17.755 1.610 ;
        RECT 14.605 0.810 17.095 1.040 ;
        RECT 20.585 0.800 20.815 1.985 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4
MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.760 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 2.430 3.210 2.710 ;
        RECT 2.950 2.200 4.075 2.430 ;
        RECT 2.950 1.770 3.210 2.200 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.898000 ;
    PORT
      LAYER Metal1 ;
        RECT 21.430 1.770 21.795 2.710 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.145 0.940 2.710 ;
        RECT 0.150 1.770 0.410 2.145 ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.745 1.770 20.010 2.710 ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.770 2.090 2.710 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.310 2.330 7.130 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 24.775 2.560 25.050 4.075 ;
        RECT 24.775 2.330 25.515 2.560 ;
        RECT 25.285 0.845 25.515 2.330 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 25.760 5.490 ;
        RECT 1.340 3.435 1.570 4.590 ;
        RECT 5.110 3.905 5.340 4.590 ;
        RECT 7.030 4.005 7.370 4.590 ;
        RECT 12.125 4.330 12.355 4.590 ;
        RECT 15.245 4.505 15.475 4.590 ;
        RECT 19.275 4.070 19.505 4.590 ;
        RECT 21.480 4.265 21.820 4.590 ;
        RECT 23.575 3.740 23.805 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 26.190 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 26.190 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.335 0.450 1.675 1.080 ;
        RECT 5.530 0.450 5.760 0.535 ;
        RECT 7.385 0.450 7.615 1.135 ;
        RECT 13.425 0.450 13.655 1.425 ;
        RECT 20.970 0.450 21.310 1.080 ;
        RECT 24.165 0.450 24.395 1.600 ;
        RECT 0.000 -0.450 25.760 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.320 3.170 0.550 4.075 ;
        RECT 3.350 3.665 3.580 4.245 ;
        RECT 10.390 4.100 10.730 4.350 ;
        RECT 15.650 4.275 17.210 4.355 ;
        RECT 15.420 4.125 17.210 4.275 ;
        RECT 19.735 4.215 20.695 4.230 ;
        RECT 15.420 4.100 15.825 4.125 ;
        RECT 5.530 3.665 9.075 3.775 ;
        RECT 3.350 3.545 9.075 3.665 ;
        RECT 3.350 3.435 5.730 3.545 ;
        RECT 0.320 2.940 4.960 3.170 ;
        RECT 6.065 2.940 7.755 3.280 ;
        RECT 2.490 1.540 2.720 2.940 ;
        RECT 4.730 2.145 4.960 2.940 ;
        RECT 7.525 2.055 7.755 2.940 ;
        RECT 8.105 2.485 8.335 3.270 ;
        RECT 8.845 2.965 9.075 3.545 ;
        RECT 9.865 3.125 10.095 3.945 ;
        RECT 10.390 3.870 15.825 4.100 ;
        RECT 19.735 4.000 21.255 4.215 ;
        RECT 10.885 3.265 13.555 3.605 ;
        RECT 14.045 3.265 15.175 3.605 ;
        RECT 9.865 2.945 10.570 3.125 ;
        RECT 9.865 2.895 14.715 2.945 ;
        RECT 10.345 2.715 14.715 2.895 ;
        RECT 8.105 2.255 9.515 2.485 ;
        RECT 0.270 1.310 2.720 1.540 ;
        RECT 6.265 1.825 7.755 2.055 ;
        RECT 8.505 2.145 9.515 2.255 ;
        RECT 0.270 0.795 0.500 1.310 ;
        RECT 6.265 1.225 6.495 1.825 ;
        RECT 6.725 1.365 8.275 1.595 ;
        RECT 3.350 0.995 3.580 1.135 ;
        RECT 6.725 0.995 6.955 1.365 ;
        RECT 3.350 0.765 6.955 0.995 ;
        RECT 8.045 0.995 8.275 1.365 ;
        RECT 8.505 1.225 8.735 2.145 ;
        RECT 9.225 0.995 9.455 1.425 ;
        RECT 10.345 1.085 10.575 2.715 ;
        RECT 14.485 2.605 14.715 2.715 ;
        RECT 10.925 1.885 11.155 2.485 ;
        RECT 11.865 2.375 12.095 2.485 ;
        RECT 14.945 2.375 15.175 3.265 ;
        RECT 11.865 2.145 16.135 2.375 ;
        RECT 10.925 1.655 15.675 1.885 ;
        RECT 8.045 0.765 9.455 0.995 ;
        RECT 15.445 0.910 15.675 1.655 ;
        RECT 15.905 1.545 16.135 2.145 ;
        RECT 16.485 1.545 16.715 3.895 ;
        RECT 17.505 3.840 17.735 3.950 ;
        RECT 19.735 3.840 19.965 4.000 ;
        RECT 20.610 3.990 21.255 4.000 ;
        RECT 20.610 3.985 23.245 3.990 ;
        RECT 17.505 3.610 19.965 3.840 ;
        RECT 17.505 1.655 17.735 3.610 ;
        RECT 18.525 2.945 18.755 3.310 ;
        RECT 15.905 1.315 16.715 1.545 ;
        RECT 17.025 1.315 17.735 1.655 ;
        RECT 18.145 2.715 19.295 2.945 ;
        RECT 18.145 1.315 18.375 2.715 ;
        RECT 18.605 0.910 18.835 2.485 ;
        RECT 15.445 0.680 18.835 0.910 ;
        RECT 19.065 1.540 19.295 2.715 ;
        RECT 20.295 1.540 20.525 3.770 ;
        RECT 21.025 3.760 23.245 3.985 ;
        RECT 19.065 1.310 20.525 1.540 ;
        RECT 20.820 1.540 21.160 2.430 ;
        RECT 22.555 1.540 22.785 3.530 ;
        RECT 23.015 2.145 23.245 3.760 ;
        RECT 24.195 2.060 24.425 2.485 ;
        RECT 23.460 1.830 24.425 2.060 ;
        RECT 23.460 1.540 23.690 1.830 ;
        RECT 20.820 1.310 23.690 1.540 ;
        RECT 19.065 0.795 19.295 1.310 ;
        RECT 23.445 0.795 23.690 1.310 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1
MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.880 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 1.770 4.330 2.290 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.123000 ;
    PORT
      LAYER Metal1 ;
        RECT 21.430 2.355 21.690 2.710 ;
        RECT 21.430 2.015 21.935 2.355 ;
        RECT 21.430 1.770 21.690 2.015 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 1.770 0.970 2.300 ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.750 1.770 20.040 2.710 ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 1.770 2.090 2.345 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.310 2.330 7.130 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 25.145 2.710 25.375 4.080 ;
        RECT 25.145 0.790 25.610 2.710 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 26.880 5.490 ;
        RECT 1.415 3.270 1.645 4.590 ;
        RECT 5.085 3.440 5.315 4.590 ;
        RECT 7.190 4.125 7.530 4.590 ;
        RECT 12.210 4.565 12.550 4.590 ;
        RECT 15.350 4.565 15.690 4.590 ;
        RECT 19.395 3.910 19.625 4.590 ;
        RECT 21.665 4.300 21.895 4.590 ;
        RECT 23.725 3.270 23.955 4.590 ;
        RECT 26.165 3.270 26.395 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.320 27.310 5.470 ;
        RECT -0.430 2.265 0.430 2.320 ;
        RECT 21.385 2.265 27.310 2.320 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 9.180 2.280 18.695 2.320 ;
        RECT 8.440 2.265 18.695 2.280 ;
        RECT -0.430 -0.430 27.310 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.075 ;
        RECT 5.505 0.450 5.735 1.080 ;
        RECT 7.545 0.450 7.775 1.080 ;
        RECT 13.545 0.450 13.775 1.480 ;
        RECT 20.970 0.450 21.310 1.080 ;
        RECT 24.165 0.450 24.395 1.600 ;
        RECT 26.405 0.450 26.635 1.600 ;
        RECT 0.000 -0.450 26.880 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 10.530 4.105 17.310 4.335 ;
        RECT 0.395 2.805 0.625 4.080 ;
        RECT 3.325 3.210 3.555 4.080 ;
        RECT 5.545 3.665 9.215 3.895 ;
        RECT 5.545 3.210 5.775 3.665 ;
        RECT 3.325 2.980 5.775 3.210 ;
        RECT 6.225 3.095 7.590 3.435 ;
        RECT 0.395 2.750 2.745 2.805 ;
        RECT 0.395 2.575 4.835 2.750 ;
        RECT 2.595 2.520 4.835 2.575 ;
        RECT 2.595 1.540 2.825 2.520 ;
        RECT 4.605 2.015 4.835 2.520 ;
        RECT 7.360 2.110 7.590 3.095 ;
        RECT 8.265 2.565 8.495 3.435 ;
        RECT 8.985 3.085 9.215 3.665 ;
        RECT 10.005 2.970 10.235 3.930 ;
        RECT 14.165 3.645 16.815 3.875 ;
        RECT 19.855 3.840 23.375 4.070 ;
        RECT 11.025 3.270 13.675 3.610 ;
        RECT 14.165 3.535 16.135 3.645 ;
        RECT 14.305 2.970 14.535 3.080 ;
        RECT 10.005 2.740 14.535 2.970 ;
        RECT 8.265 2.335 9.655 2.565 ;
        RECT 8.665 2.225 9.655 2.335 ;
        RECT 7.360 2.000 8.215 2.110 ;
        RECT 6.425 1.770 8.215 2.000 ;
        RECT 0.245 1.310 2.825 1.540 ;
        RECT 3.325 1.310 6.195 1.540 ;
        RECT 0.245 0.790 0.475 1.310 ;
        RECT 3.325 0.790 3.555 1.310 ;
        RECT 5.965 0.940 6.195 1.310 ;
        RECT 6.425 1.170 6.655 1.770 ;
        RECT 6.885 1.310 8.435 1.540 ;
        RECT 6.885 0.940 7.115 1.310 ;
        RECT 5.965 0.710 7.115 0.940 ;
        RECT 8.205 0.940 8.435 1.310 ;
        RECT 8.665 1.170 8.895 2.225 ;
        RECT 9.465 0.940 9.695 1.480 ;
        RECT 10.585 1.370 10.815 2.740 ;
        RECT 15.905 2.510 16.135 3.535 ;
        RECT 16.585 3.065 16.815 3.645 ;
        RECT 17.605 3.680 19.215 3.765 ;
        RECT 19.855 3.680 20.085 3.840 ;
        RECT 17.605 3.535 20.085 3.680 ;
        RECT 17.605 2.970 17.835 3.535 ;
        RECT 19.035 3.450 20.085 3.535 ;
        RECT 11.165 1.940 11.395 2.355 ;
        RECT 12.005 2.170 16.135 2.510 ;
        RECT 11.165 1.710 15.675 1.940 ;
        RECT 8.205 0.710 9.695 0.940 ;
        RECT 15.445 1.020 15.675 1.710 ;
        RECT 15.905 1.370 16.135 2.170 ;
        RECT 17.025 2.740 17.835 2.970 ;
        RECT 18.625 2.815 18.855 3.305 ;
        RECT 20.400 3.270 20.645 3.610 ;
        RECT 17.025 1.370 17.255 2.740 ;
        RECT 18.145 2.585 19.295 2.815 ;
        RECT 18.145 1.370 18.375 2.585 ;
        RECT 18.605 1.020 18.835 2.355 ;
        RECT 19.065 1.540 19.295 2.585 ;
        RECT 20.400 1.540 20.630 3.270 ;
        RECT 19.065 1.310 20.630 1.540 ;
        RECT 20.860 1.540 21.200 2.300 ;
        RECT 22.685 1.540 22.915 3.610 ;
        RECT 23.145 2.415 23.375 3.840 ;
        RECT 24.605 2.195 24.835 2.355 ;
        RECT 23.445 1.965 24.835 2.195 ;
        RECT 23.445 1.540 23.675 1.965 ;
        RECT 20.860 1.310 23.675 1.540 ;
        RECT 19.065 1.025 19.295 1.310 ;
        RECT 15.445 0.680 18.835 1.020 ;
        RECT 23.445 0.845 23.675 1.310 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2
MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 29.120 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 1.770 3.770 2.710 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.123000 ;
    PORT
      LAYER Metal1 ;
        RECT 21.430 2.215 21.690 3.270 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.270 0.970 2.710 ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.130 2.950 20.010 3.270 ;
        RECT 19.655 2.740 20.010 2.950 ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 2.270 2.090 2.710 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 2.890 6.570 3.270 ;
        RECT 6.280 2.530 6.570 2.890 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 24.850 3.120 25.080 4.250 ;
        RECT 26.470 3.440 27.120 4.250 ;
        RECT 26.470 3.120 26.730 3.440 ;
        RECT 24.850 2.890 27.720 3.120 ;
        RECT 25.250 0.845 25.480 2.890 ;
        RECT 27.490 0.845 27.720 2.890 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 29.120 5.490 ;
        RECT 1.265 3.440 1.495 4.590 ;
        RECT 4.950 4.560 5.290 4.590 ;
        RECT 6.885 4.560 7.225 4.590 ;
        RECT 12.120 4.510 12.350 4.590 ;
        RECT 15.320 4.510 15.550 4.590 ;
        RECT 19.390 3.985 19.620 4.590 ;
        RECT 21.595 4.375 21.935 4.590 ;
        RECT 23.710 3.440 23.940 4.590 ;
        RECT 25.870 3.440 26.100 4.590 ;
        RECT 27.910 3.440 28.140 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 29.550 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 29.550 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.535 ;
        RECT 5.445 0.450 5.675 0.530 ;
        RECT 7.460 0.450 7.690 1.380 ;
        RECT 13.460 0.450 13.690 1.535 ;
        RECT 20.990 0.450 21.220 1.255 ;
        RECT 24.130 0.450 24.360 1.525 ;
        RECT 26.370 0.450 26.600 1.650 ;
        RECT 28.610 0.450 28.840 1.650 ;
        RECT 0.000 -0.450 29.120 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.170 0.475 4.250 ;
        RECT 3.025 4.100 9.130 4.330 ;
        RECT 3.025 3.440 3.255 4.100 ;
        RECT 5.700 3.500 7.830 3.840 ;
        RECT 0.245 2.940 4.835 3.170 ;
        RECT 2.445 2.040 2.675 2.940 ;
        RECT 4.605 2.215 4.835 2.940 ;
        RECT 7.600 2.300 7.830 3.500 ;
        RECT 8.180 2.555 8.410 3.870 ;
        RECT 8.900 3.065 9.130 4.100 ;
        RECT 10.445 4.050 17.355 4.280 ;
        RECT 19.850 3.915 23.360 4.145 ;
        RECT 9.920 3.215 10.150 3.875 ;
        RECT 10.940 3.440 13.590 3.780 ;
        RECT 14.080 3.550 16.860 3.780 ;
        RECT 19.850 3.755 20.080 3.915 ;
        RECT 14.080 3.440 14.310 3.550 ;
        RECT 15.640 3.440 16.860 3.550 ;
        RECT 17.650 3.525 20.080 3.755 ;
        RECT 9.920 3.210 10.550 3.215 ;
        RECT 14.520 3.210 14.750 3.320 ;
        RECT 9.920 2.985 14.750 3.210 ;
        RECT 10.500 2.980 14.750 2.985 ;
        RECT 8.180 2.325 9.570 2.555 ;
        RECT 0.245 1.810 2.675 2.040 ;
        RECT 6.340 2.070 7.830 2.300 ;
        RECT 8.580 2.215 9.570 2.325 ;
        RECT 0.245 1.195 0.475 1.810 ;
        RECT 3.325 0.990 3.555 1.535 ;
        RECT 6.340 1.220 6.570 2.070 ;
        RECT 6.800 1.610 8.350 1.840 ;
        RECT 6.800 0.990 7.030 1.610 ;
        RECT 3.325 0.760 7.030 0.990 ;
        RECT 8.120 0.990 8.350 1.610 ;
        RECT 8.580 1.220 8.810 2.215 ;
        RECT 9.380 0.990 9.610 1.535 ;
        RECT 10.500 1.195 10.730 2.980 ;
        RECT 15.640 2.565 15.870 3.440 ;
        RECT 17.650 3.175 17.880 3.525 ;
        RECT 11.920 2.225 15.870 2.565 ;
        RECT 11.080 1.995 11.310 2.115 ;
        RECT 11.080 1.765 15.410 1.995 ;
        RECT 8.120 0.760 9.610 0.990 ;
        RECT 15.180 0.910 15.410 1.765 ;
        RECT 15.640 1.195 15.870 2.225 ;
        RECT 16.760 2.945 17.880 3.175 ;
        RECT 16.760 1.195 16.990 2.945 ;
        RECT 18.670 2.680 18.900 3.295 ;
        RECT 17.880 2.510 19.255 2.680 ;
        RECT 20.410 2.510 20.640 3.685 ;
        RECT 17.880 2.450 20.640 2.510 ;
        RECT 17.880 1.195 18.110 2.450 ;
        RECT 19.030 2.280 20.640 2.450 ;
        RECT 18.340 0.910 18.680 2.220 ;
        RECT 19.030 1.145 19.260 2.280 ;
        RECT 20.795 1.985 21.135 2.110 ;
        RECT 22.670 1.985 22.900 3.685 ;
        RECT 23.130 2.215 23.360 3.915 ;
        RECT 24.570 1.985 24.800 2.555 ;
        RECT 20.795 1.755 24.800 1.985 ;
        RECT 15.180 0.680 18.680 0.910 ;
        RECT 23.410 0.845 23.640 1.755 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4
MACRO gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.640 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 1.770 3.995 2.710 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 2.275 0.970 2.710 ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 18.630 1.770 19.425 2.710 ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 2.275 2.090 2.710 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.310 2.275 7.130 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386000 ;
    PORT
      LAYER Metal1 ;
        RECT 23.670 0.845 24.285 4.060 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 24.640 5.490 ;
        RECT 1.315 3.400 1.545 4.590 ;
        RECT 5.145 3.250 5.375 4.590 ;
        RECT 7.450 3.970 7.790 4.590 ;
        RECT 12.595 3.835 12.825 4.590 ;
        RECT 14.955 3.090 15.185 4.590 ;
        RECT 18.955 3.400 19.185 4.590 ;
        RECT 21.195 4.310 21.425 4.590 ;
        RECT 22.985 3.250 23.215 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 25.070 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 25.070 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.450 1.595 1.450 ;
        RECT 5.455 0.450 5.685 0.630 ;
        RECT 7.555 0.450 7.785 1.140 ;
        RECT 12.640 0.450 12.980 0.625 ;
        RECT 20.875 0.450 21.105 0.610 ;
        RECT 22.935 0.450 23.165 1.165 ;
        RECT 0.000 -0.450 24.640 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.295 3.170 0.525 4.060 ;
        RECT 3.325 3.630 3.555 4.210 ;
        RECT 3.325 3.400 4.915 3.630 ;
        RECT 0.295 2.940 4.455 3.170 ;
        RECT 2.545 2.045 2.775 2.940 ;
        RECT 0.245 1.815 2.775 2.045 ;
        RECT 4.225 2.070 4.455 2.940 ;
        RECT 4.685 3.020 4.915 3.400 ;
        RECT 5.605 3.510 9.675 3.740 ;
        RECT 5.605 3.020 5.835 3.510 ;
        RECT 4.685 2.790 5.835 3.020 ;
        RECT 6.485 2.940 7.675 3.280 ;
        RECT 7.445 2.505 7.675 2.940 ;
        RECT 8.575 2.505 8.805 3.235 ;
        RECT 9.445 2.930 9.675 3.510 ;
        RECT 7.445 2.275 8.280 2.505 ;
        RECT 8.575 2.275 10.170 2.505 ;
        RECT 10.515 2.285 10.745 3.730 ;
        RECT 11.095 3.605 11.325 4.360 ;
        RECT 15.735 4.020 16.865 4.360 ;
        RECT 13.025 3.605 14.725 3.720 ;
        RECT 11.095 3.490 14.725 3.605 ;
        RECT 11.095 3.375 13.225 3.490 ;
        RECT 13.935 2.745 14.165 3.260 ;
        RECT 11.880 2.515 14.165 2.745 ;
        RECT 14.495 2.860 14.725 3.490 ;
        RECT 15.735 2.860 15.965 4.020 ;
        RECT 14.495 2.630 15.965 2.860 ;
        RECT 0.245 1.110 0.475 1.815 ;
        RECT 4.225 1.730 4.835 2.070 ;
        RECT 7.445 2.060 7.675 2.275 ;
        RECT 7.215 2.045 7.675 2.060 ;
        RECT 6.435 1.830 7.675 2.045 ;
        RECT 6.435 1.815 7.300 1.830 ;
        RECT 3.325 1.090 3.555 1.450 ;
        RECT 6.435 1.140 6.665 1.815 ;
        RECT 7.385 1.585 8.245 1.600 ;
        RECT 6.895 1.370 8.245 1.585 ;
        RECT 6.895 1.355 7.470 1.370 ;
        RECT 3.325 0.910 6.210 1.090 ;
        RECT 6.895 0.910 7.125 1.355 ;
        RECT 3.325 0.860 7.125 0.910 ;
        RECT 5.985 0.680 7.125 0.860 ;
        RECT 8.015 0.910 8.245 1.370 ;
        RECT 8.575 1.140 8.905 2.275 ;
        RECT 10.515 2.055 13.640 2.285 ;
        RECT 9.395 0.910 9.625 1.135 ;
        RECT 10.515 1.025 10.745 2.055 ;
        RECT 11.195 1.085 11.425 1.825 ;
        RECT 13.935 1.545 14.165 2.515 ;
        RECT 16.195 1.910 16.425 3.730 ;
        RECT 17.215 1.940 17.445 3.900 ;
        RECT 15.055 1.680 16.425 1.910 ;
        RECT 16.835 1.710 17.445 1.940 ;
        RECT 18.170 3.170 18.465 3.900 ;
        RECT 19.975 3.170 20.205 3.950 ;
        RECT 18.170 2.940 20.205 3.170 ;
        RECT 22.215 3.020 22.445 4.100 ;
        RECT 15.055 1.545 15.285 1.680 ;
        RECT 13.935 1.315 15.285 1.545 ;
        RECT 8.015 0.680 9.625 0.910 ;
        RECT 11.195 0.855 15.780 1.085 ;
        RECT 15.440 0.680 15.780 0.855 ;
        RECT 16.175 0.910 16.405 1.450 ;
        RECT 16.835 0.910 17.065 1.710 ;
        RECT 18.170 1.480 18.400 2.940 ;
        RECT 20.555 2.790 22.445 3.020 ;
        RECT 20.555 2.220 20.785 2.790 ;
        RECT 22.215 2.560 22.445 2.790 ;
        RECT 17.295 1.140 18.985 1.480 ;
        RECT 21.635 1.070 21.865 2.560 ;
        RECT 22.215 2.220 23.440 2.560 ;
        RECT 22.215 1.110 22.445 2.220 ;
        RECT 19.205 0.910 21.865 1.070 ;
        RECT 16.175 0.840 21.865 0.910 ;
        RECT 16.175 0.680 19.425 0.840 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1
MACRO gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.200 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 1.770 4.070 2.710 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.320 1.530 2.710 ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 18.630 2.265 19.110 2.605 ;
        RECT 18.630 1.210 18.890 2.265 ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.320 2.650 2.710 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.865 2.320 7.690 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 23.605 0.845 23.930 4.050 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 25.200 5.490 ;
        RECT 1.440 3.400 1.670 4.590 ;
        RECT 5.160 3.760 5.390 4.590 ;
        RECT 7.360 3.860 7.590 4.590 ;
        RECT 12.280 3.560 12.510 4.590 ;
        RECT 14.540 3.560 14.770 4.590 ;
        RECT 18.440 3.295 18.670 4.590 ;
        RECT 20.480 3.240 20.710 4.590 ;
        RECT 22.585 3.240 22.815 4.590 ;
        RECT 24.625 3.240 24.855 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 25.630 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 25.630 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.440 0.450 1.670 1.480 ;
        RECT 5.545 0.450 5.775 0.575 ;
        RECT 7.360 0.450 7.590 1.170 ;
        RECT 12.280 0.450 12.510 1.220 ;
        RECT 20.380 0.450 20.610 1.480 ;
        RECT 22.485 0.450 22.715 1.165 ;
        RECT 24.725 0.450 24.955 1.165 ;
        RECT 0.000 -0.450 25.200 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.420 3.170 0.650 4.050 ;
        RECT 3.400 3.630 3.630 4.210 ;
        RECT 7.820 3.915 9.480 4.145 ;
        RECT 5.605 3.630 7.220 3.675 ;
        RECT 7.820 3.630 8.050 3.915 ;
        RECT 3.400 3.530 4.970 3.630 ;
        RECT 5.605 3.530 8.050 3.630 ;
        RECT 3.400 3.445 8.050 3.530 ;
        RECT 3.400 3.400 5.820 3.445 ;
        RECT 7.080 3.400 8.050 3.445 ;
        RECT 4.780 3.300 5.820 3.400 ;
        RECT 6.340 3.170 6.570 3.215 ;
        RECT 0.420 3.070 4.590 3.170 ;
        RECT 0.420 2.940 4.910 3.070 ;
        RECT 2.880 2.090 3.110 2.940 ;
        RECT 4.400 2.840 4.910 2.940 ;
        RECT 6.340 2.940 8.150 3.170 ;
        RECT 6.340 2.875 6.570 2.940 ;
        RECT 4.680 2.265 4.910 2.840 ;
        RECT 7.920 2.090 8.150 2.940 ;
        RECT 0.320 1.860 3.110 2.090 ;
        RECT 6.240 1.860 8.150 2.090 ;
        RECT 8.380 2.550 8.610 3.685 ;
        RECT 9.250 3.090 9.480 3.915 ;
        RECT 8.380 2.320 9.975 2.550 ;
        RECT 0.320 1.140 0.550 1.860 ;
        RECT 3.400 1.035 3.630 1.480 ;
        RECT 6.240 1.260 6.470 1.860 ;
        RECT 6.700 1.400 8.050 1.630 ;
        RECT 3.400 1.030 6.190 1.035 ;
        RECT 6.700 1.030 6.930 1.400 ;
        RECT 3.400 0.805 6.930 1.030 ;
        RECT 6.140 0.800 6.930 0.805 ;
        RECT 7.820 0.910 8.050 1.400 ;
        RECT 8.380 1.140 8.710 2.320 ;
        RECT 10.320 2.315 10.550 3.730 ;
        RECT 10.900 3.330 11.130 4.360 ;
        RECT 12.740 3.960 14.310 4.190 ;
        RECT 12.740 3.330 12.970 3.960 ;
        RECT 10.900 3.100 12.970 3.330 ;
        RECT 13.520 2.745 13.750 3.730 ;
        RECT 14.080 3.330 14.310 3.960 ;
        RECT 15.200 3.975 16.330 4.315 ;
        RECT 15.200 3.330 15.430 3.975 ;
        RECT 14.080 3.100 15.430 3.330 ;
        RECT 15.660 2.745 15.890 3.685 ;
        RECT 11.785 2.515 15.890 2.745 ;
        RECT 10.320 2.285 11.670 2.315 ;
        RECT 10.320 2.085 13.225 2.285 ;
        RECT 9.200 0.910 9.430 1.220 ;
        RECT 10.320 1.110 10.550 2.085 ;
        RECT 11.555 2.055 13.225 2.085 ;
        RECT 10.845 1.825 11.185 1.855 ;
        RECT 10.845 1.595 12.970 1.825 ;
        RECT 7.820 0.680 9.430 0.910 ;
        RECT 12.740 0.910 12.970 1.595 ;
        RECT 14.540 1.140 14.770 2.515 ;
        RECT 16.680 2.115 16.910 3.845 ;
        RECT 17.720 3.065 17.950 3.845 ;
        RECT 19.460 3.065 19.690 4.050 ;
        RECT 17.720 2.835 19.690 3.065 ;
        RECT 21.680 3.010 21.910 4.050 ;
        RECT 16.320 1.885 16.910 2.115 ;
        RECT 16.320 1.480 16.550 1.885 ;
        RECT 18.170 1.655 18.400 2.835 ;
        RECT 20.040 2.780 23.255 3.010 ;
        RECT 20.040 2.265 20.270 2.780 ;
        RECT 20.500 2.320 21.385 2.550 ;
        RECT 20.500 1.940 20.730 2.320 ;
        RECT 15.660 1.140 16.550 1.480 ;
        RECT 16.780 1.315 18.400 1.655 ;
        RECT 19.120 1.710 20.730 1.940 ;
        RECT 16.320 0.980 16.550 1.140 ;
        RECT 19.120 0.980 19.350 1.710 ;
        RECT 12.740 0.680 15.265 0.910 ;
        RECT 16.320 0.750 19.350 0.980 ;
        RECT 21.680 0.845 21.910 2.780 ;
        RECT 23.025 2.265 23.255 2.780 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2
MACRO gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.440 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.510 1.770 4.330 2.215 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.150 1.770 0.970 2.215 ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 18.070 1.770 18.890 2.215 ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 1.770 2.090 2.215 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.164000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 2.330 6.910 2.710 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.559650 ;
    PORT
      LAYER Metal1 ;
        RECT 23.590 3.110 23.870 3.690 ;
        RECT 25.690 3.110 25.920 3.690 ;
        RECT 23.590 2.880 25.920 3.110 ;
        RECT 23.590 1.655 23.930 2.880 ;
        RECT 23.590 1.210 26.060 1.655 ;
        RECT 23.590 0.845 23.820 1.210 ;
        RECT 25.830 0.845 26.060 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 27.440 5.490 ;
        RECT 1.315 3.230 1.545 4.590 ;
        RECT 5.085 3.400 5.315 4.590 ;
        RECT 7.200 4.125 7.540 4.590 ;
        RECT 12.045 4.510 12.275 4.590 ;
        RECT 14.305 4.070 14.535 4.590 ;
        RECT 18.305 3.075 18.535 4.590 ;
        RECT 20.565 3.880 20.795 4.590 ;
        RECT 22.605 3.880 22.835 4.590 ;
        RECT 24.660 3.880 24.890 4.590 ;
        RECT 26.850 3.880 27.080 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 27.870 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 27.870 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.450 1.650 1.075 ;
        RECT 5.505 0.450 5.735 0.530 ;
        RECT 7.305 0.450 7.535 1.180 ;
        RECT 12.225 0.450 12.455 1.120 ;
        RECT 20.230 0.450 20.460 1.265 ;
        RECT 22.470 0.450 22.700 1.655 ;
        RECT 24.710 0.450 24.940 0.980 ;
        RECT 26.950 0.450 27.180 1.655 ;
        RECT 0.000 -0.450 27.440 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 10.590 4.050 13.975 4.280 ;
        RECT 0.295 2.685 0.525 4.040 ;
        RECT 3.325 3.170 3.555 4.040 ;
        RECT 5.545 3.665 9.275 3.895 ;
        RECT 5.545 3.170 5.775 3.665 ;
        RECT 3.325 2.940 5.775 3.170 ;
        RECT 6.235 3.095 7.370 3.435 ;
        RECT 8.275 3.095 8.655 3.435 ;
        RECT 0.295 2.455 4.835 2.685 ;
        RECT 2.545 1.540 2.775 2.455 ;
        RECT 4.605 1.930 4.835 2.455 ;
        RECT 7.140 2.215 7.370 3.095 ;
        RECT 8.425 2.215 8.655 3.095 ;
        RECT 9.045 3.065 9.275 3.665 ;
        RECT 10.065 2.215 10.295 3.875 ;
        RECT 13.745 3.840 13.975 4.050 ;
        RECT 16.005 3.840 16.235 4.360 ;
        RECT 13.285 2.675 13.515 3.770 ;
        RECT 13.745 3.610 16.235 3.840 ;
        RECT 13.745 3.095 13.975 3.610 ;
        RECT 15.545 2.675 15.775 3.380 ;
        RECT 16.005 3.095 16.235 3.610 ;
        RECT 11.330 2.445 15.775 2.675 ;
        RECT 7.140 2.100 7.980 2.215 ;
        RECT 0.245 1.310 2.775 1.540 ;
        RECT 6.185 1.870 7.980 2.100 ;
        RECT 8.425 1.985 9.720 2.215 ;
        RECT 10.065 1.985 13.170 2.215 ;
        RECT 0.245 0.925 0.475 1.310 ;
        RECT 6.185 1.270 6.415 1.870 ;
        RECT 6.645 1.410 8.195 1.640 ;
        RECT 3.325 0.990 3.555 1.130 ;
        RECT 6.645 0.990 6.875 1.410 ;
        RECT 3.325 0.760 6.875 0.990 ;
        RECT 7.965 0.990 8.195 1.410 ;
        RECT 8.425 1.220 8.655 1.985 ;
        RECT 9.145 0.990 9.375 1.120 ;
        RECT 7.965 0.760 9.375 0.990 ;
        RECT 10.065 0.925 10.495 1.985 ;
        RECT 10.790 1.525 12.915 1.755 ;
        RECT 12.685 0.910 12.915 1.525 ;
        RECT 14.405 1.315 14.635 2.445 ;
        RECT 16.565 1.960 16.795 3.900 ;
        RECT 16.185 1.730 16.795 1.960 ;
        RECT 17.585 2.845 17.815 3.900 ;
        RECT 19.325 2.845 19.555 3.715 ;
        RECT 17.585 2.615 19.555 2.845 ;
        RECT 21.585 2.785 21.815 3.690 ;
        RECT 19.905 2.760 21.815 2.785 ;
        RECT 16.185 1.425 16.415 1.730 ;
        RECT 17.585 1.500 17.815 2.615 ;
        RECT 19.905 2.445 23.275 2.760 ;
        RECT 21.350 2.420 23.275 2.445 ;
        RECT 19.120 1.985 21.055 2.215 ;
        RECT 15.525 1.085 16.415 1.425 ;
        RECT 16.645 1.160 18.320 1.500 ;
        RECT 16.185 0.930 16.415 1.085 ;
        RECT 19.120 0.930 19.350 1.985 ;
        RECT 12.685 0.680 15.130 0.910 ;
        RECT 16.185 0.700 19.350 0.930 ;
        RECT 21.350 0.845 21.580 2.420 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4
MACRO gf180mcu_fd_sc_mcu9t5v0__tieh
  CLASS core TIEHIGH ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__tieh ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 2.890 1.530 3.700 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 2.240 5.490 ;
        RECT 0.250 2.945 0.480 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 2.670 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 0.450 0.480 1.355 ;
        RECT 0.000 -0.450 2.240 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.875 1.830 1.600 2.060 ;
        RECT 1.370 1.315 1.600 1.830 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__tieh
MACRO gf180mcu_fd_sc_mcu9t5v0__tiel
  CLASS core TIELOW ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__tiel ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.290400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.215 1.210 1.595 1.590 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 2.240 5.490 ;
        RECT 0.345 2.945 0.575 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 2.670 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.355 ;
        RECT 0.000 -0.450 2.240 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 2.700 1.595 3.685 ;
        RECT 0.870 2.470 1.595 2.700 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__tiel
MACRO gf180mcu_fd_sc_mcu9t5v0__xnor2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.885 2.580 3.770 2.810 ;
        RECT 1.885 2.065 2.115 2.580 ;
        RECT 3.510 2.350 3.770 2.580 ;
        RECT 3.510 2.120 4.400 2.350 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.205 3.040 4.890 3.270 ;
        RECT 1.205 2.350 1.435 3.040 ;
        RECT 4.430 2.890 4.890 3.040 ;
        RECT 0.810 2.120 1.435 2.350 ;
        RECT 4.660 2.350 4.890 2.890 ;
        RECT 4.660 2.120 5.470 2.350 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.675 3.730 3.905 4.310 ;
        RECT 3.675 3.500 5.535 3.730 ;
        RECT 5.305 2.810 5.535 3.500 ;
        RECT 5.305 2.580 6.010 2.810 ;
        RECT 5.750 1.370 6.010 2.580 ;
        RECT 4.690 1.140 6.010 1.370 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 6.720 5.490 ;
        RECT 0.285 3.500 0.515 4.590 ;
        RECT 2.325 3.500 2.555 4.590 ;
        RECT 5.765 3.500 5.995 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.150 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.150 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.325 0.450 2.555 1.355 ;
        RECT 0.000 -0.450 6.720 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.305 3.730 1.535 4.310 ;
        RECT 0.745 3.500 1.535 3.730 ;
        RECT 0.745 2.810 0.975 3.500 ;
        RECT 0.285 2.580 0.975 2.810 ;
        RECT 0.285 1.835 0.515 2.580 ;
        RECT 2.345 2.120 3.280 2.350 ;
        RECT 2.345 1.835 2.575 2.120 ;
        RECT 0.285 1.605 2.575 1.835 ;
        RECT 0.285 1.015 0.515 1.605 ;
        RECT 3.625 0.910 3.855 1.655 ;
        RECT 3.625 0.680 6.150 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor2_1
MACRO gf180mcu_fd_sc_mcu9t5v0__xnor2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.995 2.515 4.455 2.745 ;
        RECT 1.995 2.000 2.225 2.515 ;
        RECT 4.070 1.210 4.455 2.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.535 2.975 5.475 3.205 ;
        RECT 1.535 2.285 1.765 2.975 ;
        RECT 0.870 2.055 1.765 2.285 ;
        RECT 5.190 2.135 5.475 2.975 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.665 1.590 7.895 3.775 ;
        RECT 7.430 1.210 7.895 1.590 ;
        RECT 7.665 0.680 7.895 1.210 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 9.520 5.490 ;
        RECT 2.435 3.435 2.665 4.590 ;
        RECT 6.545 3.875 6.775 4.590 ;
        RECT 8.685 2.965 8.915 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 0.965 ;
        RECT 2.485 0.450 2.715 0.965 ;
        RECT 5.825 0.450 6.055 1.310 ;
        RECT 6.545 0.450 6.775 1.310 ;
        RECT 8.785 0.450 9.015 1.435 ;
        RECT 0.000 -0.450 9.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.785 4.015 6.110 4.245 ;
        RECT 0.345 1.770 0.575 3.775 ;
        RECT 3.785 3.435 4.015 4.015 ;
        RECT 4.750 3.435 5.935 3.665 ;
        RECT 2.455 2.055 3.490 2.285 ;
        RECT 5.705 2.115 5.935 3.435 ;
        RECT 2.455 1.770 2.685 2.055 ;
        RECT 5.705 1.905 7.215 2.115 ;
        RECT 0.345 1.540 2.685 1.770 ;
        RECT 4.685 1.675 7.215 1.905 ;
        RECT 1.310 0.680 1.650 1.540 ;
        RECT 4.685 0.910 4.915 1.675 ;
        RECT 3.730 0.680 4.915 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor2_2
MACRO gf180mcu_fd_sc_mcu9t5v0__xnor2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.760 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.170500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.630 3.850 2.860 ;
        RECT 1.830 1.770 2.090 2.630 ;
        RECT 3.620 2.400 3.850 2.630 ;
        RECT 3.620 2.170 4.510 2.400 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.170500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.755 3.090 4.855 3.320 ;
        RECT 0.755 2.455 0.985 3.090 ;
        RECT 4.625 2.830 4.855 3.090 ;
        RECT 4.625 2.600 5.475 2.830 ;
        RECT 0.710 1.770 0.985 2.455 ;
        RECT 5.245 2.115 5.475 2.600 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.459000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.665 3.270 7.895 3.685 ;
        RECT 7.430 2.890 7.895 3.270 ;
        RECT 7.665 1.950 7.895 2.890 ;
        RECT 9.855 1.950 10.135 3.685 ;
        RECT 7.665 1.720 10.135 1.950 ;
        RECT 7.665 0.680 7.895 1.720 ;
        RECT 9.905 0.680 10.135 1.720 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 11.760 5.490 ;
        RECT 2.665 3.875 2.895 4.590 ;
        RECT 6.645 3.875 6.875 4.590 ;
        RECT 8.735 3.875 8.965 4.590 ;
        RECT 10.925 2.875 11.155 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 12.190 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.190 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.020 ;
        RECT 2.485 0.450 2.715 1.020 ;
        RECT 5.825 0.450 6.055 1.425 ;
        RECT 6.545 0.450 6.775 1.425 ;
        RECT 8.785 0.450 9.015 1.490 ;
        RECT 11.025 0.450 11.255 1.490 ;
        RECT 0.000 -0.450 11.760 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.785 4.130 6.110 4.360 ;
        RECT 3.785 3.550 4.015 4.130 ;
        RECT 4.750 3.550 5.935 3.780 ;
        RECT 0.250 2.875 0.525 3.215 ;
        RECT 0.250 1.540 0.480 2.875 ;
        RECT 2.320 2.170 3.390 2.400 ;
        RECT 2.320 1.540 2.550 2.170 ;
        RECT 5.705 1.885 5.935 3.550 ;
        RECT 7.085 1.885 7.315 2.455 ;
        RECT 0.250 1.310 2.550 1.540 ;
        RECT 3.785 1.655 7.315 1.885 ;
        RECT 1.365 0.680 1.595 1.310 ;
        RECT 3.785 0.680 4.015 1.655 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor2_4
MACRO gf180mcu_fd_sc_mcu9t5v0__xnor3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.880 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.995 2.330 3.900 2.710 ;
        RECT 1.995 1.815 2.225 2.330 ;
        RECT 3.670 2.100 3.900 2.330 ;
        RECT 3.670 1.870 4.510 2.100 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.300 2.940 5.475 3.170 ;
        RECT 1.300 2.150 1.530 2.940 ;
        RECT 0.870 1.770 1.530 2.150 ;
        RECT 5.245 1.815 5.475 2.940 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 8.740 2.330 10.000 2.710 ;
        RECT 8.740 2.100 8.970 2.330 ;
        RECT 8.090 1.870 8.970 2.100 ;
        RECT 9.770 2.100 10.000 2.330 ;
        RECT 9.770 1.870 10.710 2.100 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.912500 ;
    PORT
      LAYER Metal1 ;
        RECT 9.985 3.720 10.215 4.360 ;
        RECT 9.985 3.645 11.855 3.720 ;
        RECT 9.985 3.490 12.190 3.645 ;
        RECT 11.685 3.415 12.190 3.490 ;
        RECT 11.960 1.590 12.190 3.415 ;
        RECT 10.950 1.210 12.190 1.590 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 12.880 5.490 ;
        RECT 2.435 3.550 2.665 4.590 ;
        RECT 6.545 3.855 6.775 4.590 ;
        RECT 8.815 3.875 9.045 4.590 ;
        RECT 12.025 3.875 12.255 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 13.310 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.310 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.080 ;
        RECT 2.485 0.450 2.715 1.080 ;
        RECT 5.825 0.450 6.055 1.080 ;
        RECT 8.585 0.450 8.815 1.080 ;
        RECT 0.000 -0.450 12.880 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.785 4.130 6.055 4.360 ;
        RECT 0.345 1.540 0.575 3.890 ;
        RECT 3.785 3.550 4.015 4.130 ;
        RECT 4.805 3.630 5.035 3.890 ;
        RECT 5.825 3.855 6.055 4.130 ;
        RECT 7.005 3.870 8.585 4.100 ;
        RECT 4.805 3.625 5.775 3.630 ;
        RECT 7.005 3.625 7.235 3.870 ;
        RECT 4.805 3.400 7.235 3.625 ;
        RECT 5.725 3.395 7.235 3.400 ;
        RECT 5.725 2.100 5.955 3.395 ;
        RECT 2.455 1.870 3.440 2.100 ;
        RECT 5.725 1.870 7.270 2.100 ;
        RECT 2.455 1.540 2.685 1.870 ;
        RECT 5.725 1.540 5.955 1.870 ;
        RECT 7.565 1.640 7.795 3.640 ;
        RECT 8.355 3.260 8.585 3.870 ;
        RECT 8.355 3.030 11.515 3.260 ;
        RECT 11.285 2.100 11.515 3.030 ;
        RECT 9.200 1.640 9.540 2.100 ;
        RECT 11.285 1.870 11.730 2.100 ;
        RECT 0.345 1.310 2.685 1.540 ;
        RECT 3.785 1.310 5.955 1.540 ;
        RECT 6.545 1.410 9.540 1.640 ;
        RECT 1.365 0.740 1.595 1.310 ;
        RECT 3.785 0.740 4.015 1.310 ;
        RECT 6.545 1.040 6.775 1.410 ;
        RECT 9.885 0.970 10.115 1.550 ;
        RECT 9.885 0.740 12.410 0.970 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor3_1
MACRO gf180mcu_fd_sc_mcu9t5v0__xnor3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.680 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.165 1.950 2.395 2.520 ;
        RECT 4.070 2.180 4.575 2.520 ;
        RECT 4.070 1.950 4.330 2.180 ;
        RECT 2.165 1.720 4.330 1.950 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.025 3.210 5.595 3.440 ;
        RECT 1.025 2.180 1.255 3.210 ;
        RECT 5.190 2.180 5.595 3.210 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 8.310 2.770 10.490 3.000 ;
        RECT 10.230 2.540 10.490 2.770 ;
        RECT 10.230 2.310 10.930 2.540 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.772000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.015 3.385 13.245 4.360 ;
        RECT 15.155 3.385 15.385 4.360 ;
        RECT 13.015 3.155 15.385 3.385 ;
        RECT 13.915 1.945 14.145 3.155 ;
        RECT 12.965 1.715 15.435 1.945 ;
        RECT 12.965 0.845 13.290 1.715 ;
        RECT 15.205 0.845 15.435 1.715 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 15.680 5.490 ;
        RECT 2.605 3.670 2.835 4.590 ;
        RECT 8.805 3.615 9.035 4.590 ;
        RECT 14.035 3.615 14.265 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 16.110 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 16.110 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.365 0.450 0.595 1.185 ;
        RECT 2.605 0.450 2.835 1.185 ;
        RECT 5.945 0.450 6.175 1.185 ;
        RECT 6.665 0.450 6.895 1.185 ;
        RECT 9.085 0.450 9.315 1.180 ;
        RECT 12.245 0.450 12.475 1.160 ;
        RECT 14.085 0.450 14.315 1.485 ;
        RECT 0.000 -0.450 15.680 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.905 4.130 6.230 4.360 ;
        RECT 0.465 1.950 0.695 3.955 ;
        RECT 3.905 3.670 4.135 4.130 ;
        RECT 4.870 3.670 6.055 3.900 ;
        RECT 1.485 2.750 3.555 2.980 ;
        RECT 1.485 1.950 1.715 2.750 ;
        RECT 3.325 2.180 3.555 2.750 ;
        RECT 5.825 2.520 6.055 3.670 ;
        RECT 6.765 2.980 6.995 4.360 ;
        RECT 12.245 3.900 12.475 4.360 ;
        RECT 10.150 3.550 12.475 3.900 ;
        RECT 6.765 2.750 8.015 2.980 ;
        RECT 11.170 2.930 12.355 3.160 ;
        RECT 7.785 2.540 8.015 2.750 ;
        RECT 5.825 2.290 7.435 2.520 ;
        RECT 0.465 1.720 1.715 1.950 ;
        RECT 1.485 0.845 1.715 1.720 ;
        RECT 7.205 1.645 7.435 2.290 ;
        RECT 4.550 1.415 7.435 1.645 ;
        RECT 4.550 1.130 4.780 1.415 ;
        RECT 3.850 0.900 4.780 1.130 ;
        RECT 7.205 0.915 7.435 1.415 ;
        RECT 7.785 2.310 9.860 2.540 ;
        RECT 12.125 2.520 12.355 2.930 ;
        RECT 7.785 1.145 8.015 2.310 ;
        RECT 11.665 2.080 11.895 2.520 ;
        RECT 8.245 1.850 11.895 2.080 ;
        RECT 12.125 2.180 13.685 2.520 ;
        RECT 8.245 0.915 8.475 1.850 ;
        RECT 12.125 1.620 12.355 2.180 ;
        RECT 7.205 0.685 8.475 0.915 ;
        RECT 10.205 1.390 12.355 1.620 ;
        RECT 10.205 0.845 10.435 1.390 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor3_2
MACRO gf180mcu_fd_sc_mcu9t5v0__xnor3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.859500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.990 2.000 2.330 2.360 ;
        RECT 3.990 2.000 4.330 2.395 ;
        RECT 1.990 1.770 4.330 2.000 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.859500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.960 3.050 3.970 3.280 ;
        RECT 0.960 2.110 1.190 3.050 ;
        RECT 3.510 2.890 3.970 3.050 ;
        RECT 3.740 2.855 3.970 2.890 ;
        RECT 3.740 2.625 5.350 2.855 ;
        RECT 5.010 2.165 5.350 2.625 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.170500 ;
    PORT
      LAYER Metal1 ;
        RECT 8.145 2.775 10.490 3.005 ;
        RECT 10.230 2.560 10.490 2.775 ;
        RECT 10.230 2.330 10.805 2.560 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.593000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.940 3.645 13.170 4.345 ;
        RECT 12.940 3.415 14.125 3.645 ;
        RECT 13.895 2.150 14.125 3.415 ;
        RECT 15.030 2.150 15.260 4.345 ;
        RECT 13.895 2.115 15.260 2.150 ;
        RECT 17.220 2.115 17.550 4.345 ;
        RECT 13.895 2.000 17.550 2.115 ;
        RECT 12.840 1.885 17.550 2.000 ;
        RECT 12.840 1.770 15.310 1.885 ;
        RECT 12.840 0.845 13.070 1.770 ;
        RECT 15.080 0.845 15.310 1.770 ;
        RECT 17.320 0.845 17.550 1.885 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.920 5.490 ;
        RECT 2.385 3.535 2.615 4.590 ;
        RECT 8.640 3.535 8.870 4.590 ;
        RECT 13.960 3.875 14.190 4.590 ;
        RECT 16.150 3.875 16.380 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 18.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 6.500 1.185 6.730 1.480 ;
        RECT 0.245 0.450 0.475 1.185 ;
        RECT 2.485 0.450 2.715 1.185 ;
        RECT 5.415 0.845 6.730 1.185 ;
        RECT 5.415 0.450 5.645 0.845 ;
        RECT 8.960 0.450 9.190 1.165 ;
        RECT 12.120 0.450 12.350 1.165 ;
        RECT 13.960 0.450 14.190 1.165 ;
        RECT 16.200 0.450 16.430 1.655 ;
        RECT 0.000 -0.450 17.920 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.605 4.105 6.110 4.335 ;
        RECT 0.345 1.880 0.575 3.875 ;
        RECT 3.605 3.535 3.835 4.105 ;
        RECT 4.625 3.315 4.855 3.875 ;
        RECT 5.880 3.535 6.110 4.105 ;
        RECT 10.080 4.130 12.350 4.360 ;
        RECT 4.625 3.085 5.810 3.315 ;
        RECT 1.420 2.590 3.290 2.820 ;
        RECT 1.420 1.880 1.650 2.590 ;
        RECT 5.580 1.940 5.810 3.085 ;
        RECT 6.600 2.910 6.830 3.875 ;
        RECT 10.080 3.550 10.310 4.130 ;
        RECT 6.600 2.680 7.850 2.910 ;
        RECT 7.620 2.545 7.850 2.680 ;
        RECT 11.100 2.545 11.330 3.900 ;
        RECT 12.120 3.550 12.350 4.130 ;
        RECT 7.040 1.940 7.270 2.450 ;
        RECT 5.580 1.935 7.270 1.940 ;
        RECT 0.345 1.650 1.650 1.880 ;
        RECT 1.365 0.845 1.650 1.650 ;
        RECT 4.560 1.710 7.270 1.935 ;
        RECT 4.560 1.705 5.630 1.710 ;
        RECT 4.560 1.130 4.790 1.705 ;
        RECT 3.550 0.900 4.790 1.130 ;
        RECT 7.040 0.910 7.270 1.710 ;
        RECT 7.620 2.315 9.785 2.545 ;
        RECT 11.100 2.315 13.665 2.545 ;
        RECT 7.620 1.140 7.850 2.315 ;
        RECT 12.055 2.230 13.665 2.315 ;
        RECT 8.080 1.855 11.825 2.085 ;
        RECT 8.080 0.910 8.310 1.855 ;
        RECT 12.055 1.625 12.285 2.230 ;
        RECT 7.040 0.680 8.310 0.910 ;
        RECT 10.080 1.395 12.285 1.625 ;
        RECT 10.080 0.815 10.310 1.395 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor3_4
MACRO gf180mcu_fd_sc_mcu9t5v0__xor2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.640 2.330 4.115 2.710 ;
        RECT 2.640 2.135 2.870 2.330 ;
        RECT 1.940 1.905 2.870 2.135 ;
        RECT 3.885 2.190 4.115 2.330 ;
        RECT 3.885 1.850 4.455 2.190 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 2.940 4.575 3.170 ;
        RECT 0.710 1.850 1.015 2.940 ;
        RECT 4.345 2.700 4.575 2.940 ;
        RECT 4.345 2.470 5.060 2.700 ;
        RECT 4.830 2.135 5.060 2.470 ;
        RECT 4.830 1.905 5.530 2.135 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.805 3.270 5.035 3.900 ;
        RECT 4.805 3.120 5.450 3.270 ;
        RECT 4.805 3.040 5.990 3.120 ;
        RECT 5.190 2.890 5.990 3.040 ;
        RECT 5.760 1.620 5.990 2.890 ;
        RECT 3.785 1.390 5.990 1.620 ;
        RECT 3.785 0.810 4.015 1.390 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 6.720 5.490 ;
        RECT 2.435 3.400 2.665 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 7.150 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.150 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.150 ;
        RECT 2.485 0.450 2.715 1.150 ;
        RECT 5.825 0.450 6.055 1.160 ;
        RECT 0.000 -0.450 6.720 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.785 4.130 6.055 4.360 ;
        RECT 0.250 3.400 0.575 3.740 ;
        RECT 3.785 3.400 4.015 4.130 ;
        RECT 5.825 3.400 6.055 4.130 ;
        RECT 0.250 1.620 0.480 3.400 ;
        RECT 3.100 1.620 3.440 2.100 ;
        RECT 0.250 1.390 3.440 1.620 ;
        RECT 1.365 0.810 1.595 1.390 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor2_1
MACRO gf180mcu_fd_sc_mcu9t5v0__xor2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.320 2.500 4.355 2.730 ;
        RECT 2.320 2.100 2.550 2.500 ;
        RECT 1.790 1.870 2.550 2.100 ;
        RECT 4.070 1.770 4.355 2.500 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.860 2.960 5.375 3.190 ;
        RECT 1.860 2.710 2.090 2.960 ;
        RECT 1.270 2.465 2.090 2.710 ;
        RECT 0.770 2.330 2.090 2.465 ;
        RECT 0.770 2.235 1.460 2.330 ;
        RECT 5.145 2.180 5.375 2.960 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.665 1.590 7.895 4.230 ;
        RECT 7.430 1.210 7.895 1.590 ;
        RECT 7.665 0.840 7.895 1.210 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 9.520 5.490 ;
        RECT 0.245 3.585 0.475 4.590 ;
        RECT 2.285 3.585 2.515 4.590 ;
        RECT 5.725 3.880 5.955 4.590 ;
        RECT 6.645 3.585 6.875 4.590 ;
        RECT 8.685 3.585 8.915 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 9.950 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.285 0.450 2.515 1.180 ;
        RECT 6.545 0.450 6.775 1.445 ;
        RECT 8.785 0.450 9.015 1.650 ;
        RECT 0.000 -0.450 9.520 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.265 3.170 1.495 4.310 ;
        RECT 3.685 3.650 3.915 4.230 ;
        RECT 3.685 3.420 5.835 3.650 ;
        RECT 0.245 2.940 1.495 3.170 ;
        RECT 0.245 1.640 0.475 2.940 ;
        RECT 2.955 1.640 3.185 2.270 ;
        RECT 5.605 2.110 5.835 3.420 ;
        RECT 5.605 1.950 7.370 2.110 ;
        RECT 4.705 1.880 7.370 1.950 ;
        RECT 4.705 1.720 5.825 1.880 ;
        RECT 0.245 1.410 3.185 1.640 ;
        RECT 0.245 0.840 0.475 1.410 ;
        RECT 3.585 0.910 3.815 1.650 ;
        RECT 4.705 1.140 4.935 1.720 ;
        RECT 5.825 0.910 6.055 1.490 ;
        RECT 3.585 0.680 6.055 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor2_2
MACRO gf180mcu_fd_sc_mcu9t5v0__xor2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.760 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.170500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.790 2.330 4.360 2.710 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.170500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.770 2.940 4.860 3.170 ;
        RECT 0.770 2.330 1.110 2.940 ;
        RECT 4.630 2.710 4.860 2.940 ;
        RECT 4.630 2.330 5.430 2.710 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.459000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.430 3.450 7.895 4.360 ;
        RECT 7.665 2.115 7.895 3.450 ;
        RECT 9.855 2.115 10.135 4.360 ;
        RECT 7.665 1.885 10.135 2.115 ;
        RECT 7.665 0.845 7.895 1.885 ;
        RECT 9.905 0.845 10.135 1.885 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 11.760 5.490 ;
        RECT 0.245 3.860 0.475 4.590 ;
        RECT 2.285 3.860 2.515 4.590 ;
        RECT 5.725 3.860 5.955 4.590 ;
        RECT 6.645 3.860 6.875 4.590 ;
        RECT 8.735 3.860 8.965 4.590 ;
        RECT 10.925 3.860 11.155 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 12.190 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.190 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.230 0.450 2.570 1.595 ;
        RECT 6.545 0.450 6.775 1.165 ;
        RECT 8.785 0.450 9.015 1.655 ;
        RECT 11.025 0.450 11.255 1.655 ;
        RECT 0.000 -0.450 11.760 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.265 3.630 1.495 4.065 ;
        RECT 0.190 3.400 1.495 3.630 ;
        RECT 3.635 3.630 3.865 4.360 ;
        RECT 3.635 3.400 5.890 3.630 ;
        RECT 0.190 2.100 0.420 3.400 ;
        RECT 5.660 2.210 5.890 3.400 ;
        RECT 5.660 2.100 7.315 2.210 ;
        RECT 0.190 1.870 3.290 2.100 ;
        RECT 4.705 1.870 7.315 2.100 ;
        RECT 0.190 1.365 0.530 1.870 ;
        RECT 3.585 1.060 3.815 1.650 ;
        RECT 4.705 1.310 4.935 1.870 ;
        RECT 5.825 1.060 6.055 1.640 ;
        RECT 3.585 0.830 6.055 1.060 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor2_4
MACRO gf180mcu_fd_sc_mcu9t5v0__xor3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.880 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.890 1.770 2.650 2.155 ;
        RECT 2.420 1.640 2.650 1.770 ;
        RECT 4.225 1.640 4.455 2.210 ;
        RECT 2.420 1.410 4.455 1.640 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.925 3.075 1.530 3.270 ;
        RECT 0.925 2.845 5.475 3.075 ;
        RECT 0.925 1.870 1.155 2.845 ;
        RECT 5.245 1.870 5.475 2.845 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 7.990 2.480 10.755 2.710 ;
        RECT 7.990 2.330 8.335 2.480 ;
        RECT 10.525 1.870 10.755 2.480 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.105 3.270 11.335 3.700 ;
        RECT 11.105 2.890 12.235 3.270 ;
        RECT 12.005 1.155 12.235 2.890 ;
        RECT 10.030 0.925 12.235 1.155 ;
        RECT 10.030 0.895 10.370 0.925 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 12.880 5.490 ;
        RECT 2.385 3.305 2.615 4.590 ;
        RECT 8.685 2.965 8.915 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 13.310 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.310 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.180 ;
        RECT 2.485 0.450 2.715 1.180 ;
        RECT 5.825 0.450 6.055 1.180 ;
        RECT 6.545 0.450 6.775 1.180 ;
        RECT 8.785 0.450 9.015 1.180 ;
        RECT 12.125 0.450 12.355 0.695 ;
        RECT 0.000 -0.450 12.880 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.785 3.830 6.110 4.115 ;
        RECT 10.085 4.005 12.635 4.235 ;
        RECT 0.345 1.640 0.575 3.645 ;
        RECT 3.785 3.305 4.015 3.830 ;
        RECT 4.750 3.360 5.935 3.590 ;
        RECT 1.385 2.385 3.335 2.615 ;
        RECT 1.385 1.640 1.615 2.385 ;
        RECT 3.105 1.870 3.335 2.385 ;
        RECT 5.705 1.640 5.935 3.360 ;
        RECT 6.630 2.670 6.860 3.775 ;
        RECT 10.085 3.305 10.315 4.005 ;
        RECT 12.405 3.425 12.635 4.005 ;
        RECT 6.630 2.440 7.760 2.670 ;
        RECT 7.070 1.640 7.300 2.210 ;
        RECT 7.530 2.100 7.760 2.440 ;
        RECT 9.400 2.100 9.740 2.155 ;
        RECT 7.530 1.890 9.740 2.100 ;
        RECT 0.345 1.410 1.615 1.640 ;
        RECT 1.365 0.840 1.615 1.410 ;
        RECT 4.685 1.620 7.300 1.640 ;
        RECT 7.665 1.870 9.740 1.890 ;
        RECT 4.685 1.410 7.435 1.620 ;
        RECT 4.685 1.125 4.915 1.410 ;
        RECT 3.730 0.895 4.915 1.125 ;
        RECT 7.205 0.910 7.435 1.410 ;
        RECT 7.665 1.140 7.895 1.870 ;
        RECT 11.545 1.640 11.775 2.210 ;
        RECT 8.325 1.410 11.775 1.640 ;
        RECT 8.325 0.910 8.555 1.410 ;
        RECT 7.205 0.680 8.555 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor3_1
MACRO gf180mcu_fd_sc_mcu9t5v0__xor3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.680 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 1.740 2.170 2.200 ;
        RECT 4.225 1.740 4.455 2.025 ;
        RECT 1.830 1.510 4.455 1.740 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.910 2.890 3.900 3.270 ;
        RECT 0.910 1.915 1.140 2.890 ;
        RECT 3.670 2.485 3.900 2.890 ;
        RECT 3.670 2.255 5.530 2.485 ;
        RECT 5.190 1.970 5.530 2.255 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.560500 ;
    PORT
      LAYER Metal1 ;
        RECT 8.090 2.370 10.710 2.710 ;
        RECT 9.670 2.330 10.710 2.370 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.772000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.845 3.645 13.075 4.320 ;
        RECT 12.845 3.415 14.030 3.645 ;
        RECT 13.800 1.670 14.030 3.415 ;
        RECT 14.985 1.670 15.315 3.685 ;
        RECT 12.845 1.440 15.315 1.670 ;
        RECT 12.845 0.845 13.290 1.440 ;
        RECT 15.085 0.845 15.315 1.440 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 15.680 5.490 ;
        RECT 2.435 3.510 2.665 4.590 ;
        RECT 6.545 3.450 6.775 4.590 ;
        RECT 8.815 4.350 9.045 4.590 ;
        RECT 12.025 4.350 12.255 4.590 ;
        RECT 13.865 3.875 14.095 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 16.110 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 16.110 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.185 ;
        RECT 2.485 0.450 2.715 1.185 ;
        RECT 5.825 0.450 6.055 1.185 ;
        RECT 8.585 0.450 8.815 1.185 ;
        RECT 13.965 0.450 14.195 1.165 ;
        RECT 0.000 -0.450 15.680 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.785 4.130 6.055 4.360 ;
        RECT 0.345 1.685 0.575 3.850 ;
        RECT 3.785 3.510 4.015 4.130 ;
        RECT 4.805 2.945 5.035 3.900 ;
        RECT 5.825 3.175 6.055 4.130 ;
        RECT 9.930 4.135 11.360 4.155 ;
        RECT 9.930 3.925 11.940 4.135 ;
        RECT 11.265 3.905 11.940 3.925 ;
        RECT 7.005 3.465 11.170 3.695 ;
        RECT 7.005 2.945 7.235 3.465 ;
        RECT 4.805 2.715 7.235 2.945 ;
        RECT 1.370 2.430 3.440 2.660 ;
        RECT 1.370 1.685 1.600 2.430 ;
        RECT 3.100 1.970 3.440 2.430 ;
        RECT 0.345 1.455 1.600 1.685 ;
        RECT 7.005 1.645 7.235 2.715 ;
        RECT 1.365 0.845 1.600 1.455 ;
        RECT 4.685 1.415 7.235 1.645 ;
        RECT 7.565 2.140 7.795 3.235 ;
        RECT 10.940 2.410 11.170 3.465 ;
        RECT 11.710 2.870 11.940 3.905 ;
        RECT 11.710 2.640 12.190 2.870 ;
        RECT 10.940 2.180 11.730 2.410 ;
        RECT 7.565 1.910 9.540 2.140 ;
        RECT 11.960 2.130 12.190 2.640 ;
        RECT 11.960 1.950 13.570 2.130 ;
        RECT 4.685 1.130 4.915 1.415 ;
        RECT 7.565 1.130 7.795 1.910 ;
        RECT 11.005 1.900 13.570 1.950 ;
        RECT 11.005 1.720 12.185 1.900 ;
        RECT 3.730 0.900 4.915 1.130 ;
        RECT 6.490 0.900 7.795 1.130 ;
        RECT 9.885 0.910 10.115 1.655 ;
        RECT 11.005 1.140 11.235 1.720 ;
        RECT 12.125 0.910 12.355 1.490 ;
        RECT 9.885 0.680 12.355 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor3_2
MACRO gf180mcu_fd_sc_mcu9t5v0__xor3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.859500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.005 2.170 2.135 ;
        RECT 4.045 2.005 4.275 2.520 ;
        RECT 1.830 1.775 4.275 2.005 ;
        RECT 1.830 1.210 2.090 1.775 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.859500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.905 3.005 2.880 3.055 ;
        RECT 0.905 2.825 4.860 3.005 ;
        RECT 0.905 2.180 1.135 2.825 ;
        RECT 2.735 2.775 4.860 2.825 ;
        RECT 4.630 2.710 4.860 2.775 ;
        RECT 4.630 2.180 5.295 2.710 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.170500 ;
    PORT
      LAYER Metal1 ;
        RECT 7.910 2.475 10.480 2.710 ;
        RECT 9.670 2.330 10.480 2.475 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.593000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.765 3.465 12.995 4.360 ;
        RECT 12.765 3.235 13.950 3.465 ;
        RECT 13.720 2.030 13.950 3.235 ;
        RECT 14.955 2.115 15.185 4.360 ;
        RECT 17.045 2.115 17.375 4.360 ;
        RECT 14.955 2.030 17.375 2.115 ;
        RECT 13.720 1.885 17.375 2.030 ;
        RECT 13.720 1.720 15.135 1.885 ;
        RECT 13.590 1.490 15.135 1.720 ;
        RECT 12.665 1.210 15.135 1.490 ;
        RECT 12.665 0.680 12.895 1.210 ;
        RECT 14.905 0.845 15.135 1.210 ;
        RECT 17.145 0.845 17.375 1.885 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.590 17.920 5.490 ;
        RECT 2.385 3.695 2.615 4.590 ;
        RECT 6.365 3.015 6.595 4.590 ;
        RECT 8.685 3.865 8.915 4.590 ;
        RECT 11.845 4.350 12.075 4.590 ;
        RECT 13.785 3.695 14.015 4.590 ;
        RECT 15.975 3.695 16.205 4.590 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.265 18.350 5.470 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 2.265 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.450 0.475 1.185 ;
        RECT 2.485 0.450 2.715 1.185 ;
        RECT 5.645 0.450 5.875 1.185 ;
        RECT 8.405 0.450 8.635 1.185 ;
        RECT 13.785 0.450 14.015 0.695 ;
        RECT 16.025 0.450 16.255 1.655 ;
        RECT 0.000 -0.450 17.920 0.450 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.605 4.130 5.875 4.360 ;
        RECT 0.345 1.950 0.575 4.035 ;
        RECT 3.605 3.695 3.835 4.130 ;
        RECT 4.625 3.465 4.855 3.900 ;
        RECT 5.645 3.695 5.875 4.130 ;
        RECT 9.700 3.865 11.955 4.095 ;
        RECT 6.825 3.635 8.545 3.680 ;
        RECT 4.625 3.235 5.755 3.465 ;
        RECT 1.365 2.465 2.590 2.595 ;
        RECT 1.365 2.365 3.310 2.465 ;
        RECT 1.365 1.950 1.595 2.365 ;
        RECT 2.380 2.235 3.310 2.365 ;
        RECT 5.525 2.410 5.755 3.235 ;
        RECT 6.825 3.450 11.495 3.635 ;
        RECT 6.825 2.410 7.055 3.450 ;
        RECT 8.405 3.405 11.495 3.450 ;
        RECT 0.345 1.720 1.595 1.950 ;
        RECT 1.365 0.845 1.595 1.720 ;
        RECT 5.525 2.180 7.055 2.410 ;
        RECT 7.385 2.245 7.615 3.220 ;
        RECT 5.525 1.645 5.755 2.180 ;
        RECT 7.385 2.015 9.410 2.245 ;
        RECT 11.265 2.180 11.495 3.405 ;
        RECT 11.725 2.160 11.955 3.865 ;
        RECT 7.385 1.950 7.615 2.015 ;
        RECT 11.725 1.950 13.490 2.160 ;
        RECT 4.465 1.415 5.755 1.645 ;
        RECT 6.365 1.720 7.615 1.950 ;
        RECT 10.825 1.930 13.490 1.950 ;
        RECT 10.825 1.720 11.955 1.930 ;
        RECT 4.465 1.130 4.695 1.415 ;
        RECT 3.550 0.900 4.695 1.130 ;
        RECT 6.365 0.845 6.595 1.720 ;
        RECT 9.705 0.910 9.935 1.655 ;
        RECT 10.825 1.315 11.055 1.720 ;
        RECT 11.945 0.910 12.175 1.490 ;
        RECT 9.705 0.680 12.175 0.910 ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor3_4
SITE GF018hv5v_mcu_sc7
  SYMMETRY X Y ;
  CLASS core ;
  SIZE 0.56 BY 3.92 ;
END GF018hv5v_mcu_sc7
MACRO gf180mcu_fd_sc_mcu7t5v0__addf_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__addf_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.480 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.272000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.615 1.770 3.470 2.150 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.272000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.640 1.795 17.070 2.150 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.694000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.890 1.620 13.910 1.850 ;
        RECT 12.340 1.200 13.910 1.620 ;
        RECT 13.540 0.550 13.910 1.200 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.893200 ;
    PORT
      LAYER Metal1 ;
        RECT 17.450 0.790 17.830 3.370 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.847000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.140 0.610 0.575 3.370 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 18.480 4.220 ;
        RECT 1.365 3.040 1.595 3.620 ;
        RECT 6.790 3.005 7.130 3.620 ;
        RECT 9.105 2.705 9.335 3.620 ;
        RECT 11.310 3.005 11.650 3.620 ;
        RECT 16.445 2.480 16.675 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 18.910 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.910 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 0.870 ;
        RECT 6.790 0.300 7.130 0.915 ;
        RECT 9.250 0.300 9.590 1.090 ;
        RECT 11.310 0.300 11.650 0.915 ;
        RECT 16.445 0.300 16.675 0.765 ;
        RECT 0.000 -0.300 18.480 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.925 2.560 4.710 2.790 ;
        RECT 5.550 2.775 5.890 2.845 ;
        RECT 8.030 2.775 8.370 2.845 ;
        RECT 0.925 1.390 1.155 2.560 ;
        RECT 5.550 2.545 8.370 2.775 ;
        RECT 10.070 2.545 13.430 2.775 ;
        RECT 14.165 2.315 14.400 2.765 ;
        RECT 5.010 2.080 14.400 2.315 ;
        RECT 14.170 1.565 14.400 2.080 ;
        RECT 0.925 1.160 4.615 1.390 ;
        RECT 4.385 0.810 4.615 1.160 ;
        RECT 5.505 1.145 8.415 1.375 ;
        RECT 5.505 0.810 5.735 1.145 ;
        RECT 8.185 0.810 8.415 1.145 ;
        RECT 10.025 1.145 12.110 1.375 ;
        RECT 10.025 0.770 10.255 1.145 ;
        RECT 11.880 0.915 12.110 1.145 ;
        RECT 14.170 1.335 17.200 1.565 ;
        RECT 11.880 0.680 13.210 0.915 ;
        RECT 14.170 0.750 14.495 1.335 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__addf_1
MACRO gf180mcu_fd_sc_mcu7t5v0__addf_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__addf_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.160 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.372000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.605 1.760 4.130 2.160 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.372000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.340 2.160 16.700 3.370 ;
        RECT 15.580 1.760 17.335 2.160 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.754000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.490 1.835 5.660 2.160 ;
        RECT 4.490 1.605 14.755 1.835 ;
        RECT 14.525 1.345 14.755 1.605 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.045200 ;
    PORT
      LAYER Metal1 ;
        RECT 18.370 0.550 18.960 3.370 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.006200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.220 0.550 1.680 3.370 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 20.160 4.220 ;
        RECT 0.385 2.460 0.615 3.620 ;
        RECT 2.370 3.285 2.710 3.620 ;
        RECT 7.950 3.005 8.290 3.620 ;
        RECT 10.530 2.845 10.870 3.620 ;
        RECT 12.490 3.005 12.830 3.620 ;
        RECT 17.405 2.480 17.635 3.620 ;
        RECT 19.445 2.480 19.675 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 20.590 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 20.590 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.285 0.300 0.515 0.905 ;
        RECT 2.525 0.300 2.755 0.695 ;
        RECT 7.950 0.300 8.290 0.915 ;
        RECT 10.530 0.300 10.870 1.075 ;
        RECT 12.590 0.300 12.930 0.915 ;
        RECT 17.230 0.300 17.570 0.730 ;
        RECT 19.545 0.300 19.775 0.905 ;
        RECT 0.000 -0.300 20.160 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.940 2.610 5.830 2.845 ;
        RECT 1.940 1.155 2.170 2.610 ;
        RECT 6.710 2.540 9.790 2.775 ;
        RECT 11.240 2.545 14.310 2.775 ;
        RECT 15.105 2.295 15.335 3.140 ;
        RECT 6.070 2.065 15.335 2.295 ;
        RECT 1.940 0.925 5.775 1.155 ;
        RECT 5.545 0.780 5.775 0.925 ;
        RECT 6.665 1.145 9.695 1.375 ;
        RECT 6.665 0.790 6.895 1.145 ;
        RECT 9.465 0.790 9.695 1.145 ;
        RECT 11.305 1.145 14.215 1.375 ;
        RECT 11.305 0.790 11.535 1.145 ;
        RECT 13.985 0.790 14.215 1.145 ;
        RECT 15.105 1.315 15.335 2.065 ;
        RECT 17.890 1.315 18.120 2.230 ;
        RECT 15.105 1.085 18.120 1.315 ;
        RECT 15.105 0.780 15.335 1.085 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__addf_2
MACRO gf180mcu_fd_sc_mcu7t5v0__addf_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__addf_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.640 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.352000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.095 1.770 6.785 2.150 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.352000 ;
    PORT
      LAYER Metal1 ;
        RECT 17.450 1.770 19.650 2.160 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.734000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.330 1.625 17.110 1.855 ;
        RECT 12.325 0.650 12.755 1.625 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.597200 ;
    PORT
      LAYER Metal1 ;
        RECT 20.790 2.240 21.260 3.370 ;
        RECT 23.030 2.240 23.410 3.370 ;
        RECT 20.790 1.920 23.410 2.240 ;
        RECT 23.030 1.135 23.410 1.920 ;
        RECT 20.805 0.905 23.410 1.135 ;
        RECT 20.805 0.530 21.035 0.905 ;
        RECT 23.030 0.530 23.410 0.905 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.424400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.215 2.240 1.675 3.370 ;
        RECT 3.460 2.240 3.915 3.370 ;
        RECT 1.215 1.920 3.915 2.240 ;
        RECT 1.215 1.135 1.675 1.920 ;
        RECT 1.215 0.905 3.915 1.135 ;
        RECT 1.215 0.530 1.675 0.905 ;
        RECT 3.685 0.530 3.915 0.905 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 24.640 4.220 ;
        RECT 0.325 2.650 0.555 3.620 ;
        RECT 2.565 2.650 2.795 3.620 ;
        RECT 4.805 3.160 5.035 3.620 ;
        RECT 10.230 3.005 10.570 3.620 ;
        RECT 12.765 2.670 12.995 3.620 ;
        RECT 14.990 3.005 15.330 3.620 ;
        RECT 19.585 3.160 19.815 3.620 ;
        RECT 21.925 2.560 22.155 3.620 ;
        RECT 24.165 2.560 24.395 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 25.070 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 25.070 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.325 0.300 0.555 0.870 ;
        RECT 2.505 0.300 2.850 0.675 ;
        RECT 4.750 0.300 5.090 0.675 ;
        RECT 10.230 0.300 10.570 0.915 ;
        RECT 12.985 0.300 13.215 1.135 ;
        RECT 14.990 0.300 15.330 0.915 ;
        RECT 19.685 0.300 19.915 0.765 ;
        RECT 21.870 0.300 22.210 0.670 ;
        RECT 24.165 0.300 24.395 0.765 ;
        RECT 0.000 -0.300 24.640 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 8.990 2.775 9.330 2.830 ;
        RECT 11.590 2.775 11.930 2.830 ;
        RECT 4.560 2.545 8.110 2.775 ;
        RECT 8.990 2.545 11.930 2.775 ;
        RECT 13.740 2.545 16.570 2.775 ;
        RECT 16.935 2.550 20.355 2.785 ;
        RECT 4.560 1.670 4.790 2.545 ;
        RECT 16.935 2.315 17.165 2.550 ;
        RECT 8.380 2.085 17.165 2.315 ;
        RECT 1.915 1.440 4.790 1.670 ;
        RECT 4.560 1.140 4.790 1.440 ;
        RECT 20.125 1.670 20.355 2.550 ;
        RECT 20.125 1.440 22.785 1.670 ;
        RECT 8.945 1.145 11.860 1.375 ;
        RECT 4.560 0.905 8.110 1.140 ;
        RECT 7.770 0.780 8.110 0.905 ;
        RECT 8.945 0.795 9.175 1.145 ;
        RECT 11.630 0.795 11.860 1.145 ;
        RECT 13.705 1.145 16.615 1.375 ;
        RECT 20.125 1.365 20.355 1.440 ;
        RECT 13.705 0.810 13.935 1.145 ;
        RECT 16.385 0.810 16.615 1.145 ;
        RECT 17.505 1.135 20.355 1.365 ;
        RECT 17.505 0.810 17.735 1.135 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__addf_4
MACRO gf180mcu_fd_sc_mcu7t5v0__addh_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__addh_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.175000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.775 2.365 6.095 2.595 ;
        RECT 2.775 2.150 3.270 2.365 ;
        RECT 1.505 1.770 3.270 2.150 ;
        RECT 5.865 1.870 6.095 2.365 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.175000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.725 1.790 5.510 2.135 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.895400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.140 0.650 0.575 3.370 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.895400 ;
    PORT
      LAYER Metal1 ;
        RECT 9.405 1.680 9.735 3.370 ;
        RECT 8.975 0.650 9.735 1.680 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 10.080 4.220 ;
        RECT 1.365 3.230 1.595 3.620 ;
        RECT 3.590 3.285 3.930 3.620 ;
        RECT 4.330 3.285 4.670 3.620 ;
        RECT 8.205 3.075 8.435 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 10.510 4.350 ;
        RECT -0.430 1.760 5.190 1.885 ;
        RECT 6.710 1.760 10.510 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 5.190 1.760 6.710 1.885 ;
        RECT -0.430 -0.430 10.510 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.640 ;
        RECT 8.150 0.300 8.490 1.035 ;
        RECT 0.000 -0.300 10.080 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.140 3.100 3.340 3.330 ;
        RECT 2.140 3.000 2.370 3.100 ;
        RECT 0.925 2.770 2.370 3.000 ;
        RECT 3.110 3.055 3.340 3.100 ;
        RECT 3.110 2.825 6.645 3.055 ;
        RECT 7.010 3.010 7.350 3.240 ;
        RECT 0.925 1.100 1.155 2.770 ;
        RECT 6.415 1.970 6.645 2.825 ;
        RECT 7.120 2.610 7.350 3.010 ;
        RECT 7.120 2.375 8.370 2.610 ;
        RECT 8.140 2.250 8.370 2.375 ;
        RECT 6.415 1.740 7.910 1.970 ;
        RECT 8.140 1.910 9.055 2.250 ;
        RECT 8.140 1.495 8.370 1.910 ;
        RECT 5.570 1.265 8.370 1.495 ;
        RECT 0.925 0.870 3.850 1.100 ;
        RECT 3.475 0.810 3.850 0.870 ;
        RECT 4.230 0.760 4.570 1.035 ;
        RECT 5.570 0.990 5.910 1.265 ;
        RECT 6.910 0.760 7.250 1.035 ;
        RECT 4.230 0.530 7.250 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__addh_1
MACRO gf180mcu_fd_sc_mcu7t5v0__addh_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__addh_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.320 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.073000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.435 2.350 7.770 2.710 ;
        RECT 3.435 2.150 3.780 2.350 ;
        RECT 7.380 2.205 7.770 2.350 ;
        RECT 2.715 1.740 3.780 2.150 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.073000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.010 1.720 5.620 2.120 ;
        RECT 4.010 1.210 4.390 1.720 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.177100 ;
    PORT
      LAYER Metal1 ;
        RECT 1.210 0.550 1.615 3.370 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.930800 ;
    PORT
      LAYER Metal1 ;
        RECT 10.490 2.480 11.110 3.370 ;
        RECT 10.490 2.250 11.650 2.480 ;
        RECT 11.310 1.560 11.650 2.250 ;
        RECT 10.490 1.220 11.650 1.560 ;
        RECT 10.490 0.550 11.110 1.220 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 12.320 4.220 ;
        RECT 0.315 2.480 0.545 3.620 ;
        RECT 2.400 3.215 2.740 3.620 ;
        RECT 4.490 3.215 4.830 3.620 ;
        RECT 5.430 3.215 5.770 3.620 ;
        RECT 9.370 2.685 9.710 3.620 ;
        RECT 11.510 2.710 11.850 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 12.750 4.350 ;
        RECT -0.430 1.760 6.200 1.885 ;
        RECT 7.425 1.760 12.750 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 6.200 1.760 7.425 1.885 ;
        RECT -0.430 -0.430 12.750 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.265 0.300 0.495 0.985 ;
        RECT 2.505 0.300 2.735 0.940 ;
        RECT 9.425 0.300 9.655 0.780 ;
        RECT 11.665 0.300 11.895 0.780 ;
        RECT 0.000 -0.300 12.320 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.975 2.985 3.810 3.170 ;
        RECT 2.015 2.940 3.810 2.985 ;
        RECT 2.015 2.755 3.205 2.940 ;
        RECT 2.015 1.410 2.245 2.755 ;
        RECT 8.010 2.435 8.350 3.370 ;
        RECT 8.010 2.205 9.400 2.435 ;
        RECT 9.170 2.020 9.400 2.205 ;
        RECT 6.095 1.745 8.790 1.975 ;
        RECT 9.170 1.790 10.790 2.020 ;
        RECT 6.095 1.420 6.325 1.745 ;
        RECT 9.170 1.515 9.400 1.790 ;
        RECT 2.015 1.180 3.355 1.410 ;
        RECT 3.125 0.760 3.355 1.180 ;
        RECT 4.665 1.190 6.325 1.420 ;
        RECT 6.670 1.285 9.400 1.515 ;
        RECT 4.665 0.760 4.895 1.190 ;
        RECT 6.670 0.990 7.010 1.285 ;
        RECT 3.125 0.530 4.895 0.760 ;
        RECT 5.330 0.530 8.350 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__addh_2
MACRO gf180mcu_fd_sc_mcu7t5v0__addh_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__addh_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.400 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.696000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 2.015 10.470 2.245 ;
        RECT 1.100 1.685 1.330 2.015 ;
        RECT 3.905 1.800 5.845 2.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.696000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.640 1.570 3.470 1.775 ;
        RECT 6.355 1.570 7.620 1.785 ;
        RECT 1.640 1.555 7.620 1.570 ;
        RECT 1.640 1.305 6.585 1.555 ;
        RECT 1.640 1.200 3.965 1.305 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.270100 ;
    PORT
      LAYER Metal1 ;
        RECT 13.170 2.150 13.510 2.885 ;
        RECT 15.850 2.150 16.240 2.885 ;
        RECT 13.170 1.770 16.240 2.150 ;
        RECT 13.170 1.035 13.560 1.770 ;
        RECT 15.900 1.035 16.240 1.770 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.090300 ;
    PORT
      LAYER Metal1 ;
        RECT 18.220 2.480 18.560 3.390 ;
        RECT 20.250 2.480 20.845 3.390 ;
        RECT 18.220 2.245 20.845 2.480 ;
        RECT 20.250 1.370 20.845 2.245 ;
        RECT 18.220 1.135 20.845 1.370 ;
        RECT 18.220 0.540 18.605 1.135 ;
        RECT 20.250 0.650 20.845 1.135 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 22.400 4.220 ;
        RECT 0.245 3.145 0.475 3.620 ;
        RECT 2.335 3.105 2.565 3.620 ;
        RECT 4.425 3.105 4.655 3.620 ;
        RECT 8.300 3.445 8.640 3.620 ;
        RECT 12.045 3.285 12.385 3.620 ;
        RECT 14.510 3.285 14.850 3.620 ;
        RECT 17.125 2.730 17.355 3.620 ;
        RECT 19.395 2.730 19.625 3.620 ;
        RECT 21.605 2.730 21.835 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.990 22.830 4.350 ;
        RECT -0.430 1.760 3.980 1.990 ;
        RECT 17.930 1.760 22.830 1.990 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 3.980 1.760 17.930 1.990 ;
        RECT -0.430 -0.430 22.830 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 0.690 ;
        RECT 4.370 0.300 4.710 1.075 ;
        RECT 12.090 0.300 12.440 1.120 ;
        RECT 14.560 0.300 14.900 0.635 ;
        RECT 17.225 0.300 17.455 0.935 ;
        RECT 19.440 0.300 19.780 0.735 ;
        RECT 21.735 0.300 21.965 0.935 ;
        RECT 0.000 -0.300 22.400 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.255 2.815 1.600 3.390 ;
        RECT 3.350 2.815 3.690 3.390 ;
        RECT 5.720 3.055 11.615 3.215 ;
        RECT 12.660 3.115 14.055 3.345 ;
        RECT 12.660 3.055 12.890 3.115 ;
        RECT 5.720 2.985 12.890 3.055 ;
        RECT 11.385 2.825 12.890 2.985 ;
        RECT 13.825 2.980 14.055 3.115 ;
        RECT 15.315 3.115 16.700 3.345 ;
        RECT 15.315 2.980 15.545 3.115 ;
        RECT 0.640 2.755 3.690 2.815 ;
        RECT 0.640 2.525 10.930 2.755 ;
        RECT 13.825 2.750 15.545 2.980 ;
        RECT 0.640 1.320 0.870 2.525 ;
        RECT 10.700 2.045 10.930 2.525 ;
        RECT 10.700 1.815 12.880 2.045 ;
        RECT 16.470 1.970 16.700 3.115 ;
        RECT 16.470 1.740 19.860 1.970 ;
        RECT 9.640 1.380 12.920 1.585 ;
        RECT 7.885 1.350 12.920 1.380 ;
        RECT 7.885 1.325 9.980 1.350 ;
        RECT 0.640 1.090 1.255 1.320 ;
        RECT 6.840 1.145 9.980 1.325 ;
        RECT 6.840 1.090 8.115 1.145 ;
        RECT 9.640 1.090 9.980 1.145 ;
        RECT 1.025 0.770 1.255 1.090 ;
        RECT 5.720 0.860 6.060 1.075 ;
        RECT 8.300 0.860 8.640 0.915 ;
        RECT 10.760 0.860 11.100 1.075 ;
        RECT 1.025 0.540 2.670 0.770 ;
        RECT 5.720 0.630 11.100 0.860 ;
        RECT 12.690 0.760 12.920 1.350 ;
        RECT 14.030 1.005 15.565 1.235 ;
        RECT 14.030 0.760 14.260 1.005 ;
        RECT 12.690 0.530 14.260 0.760 ;
        RECT 15.335 0.760 15.565 1.005 ;
        RECT 16.470 0.760 16.700 1.740 ;
        RECT 15.335 0.530 16.700 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__addh_4
MACRO gf180mcu_fd_sc_mcu7t5v0__and2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.519000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.660 1.540 1.020 2.810 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.519000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.780 1.540 2.140 3.370 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.893200 ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 0.555 3.870 3.380 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 4.480 4.220 ;
        RECT 0.245 3.225 0.475 3.620 ;
        RECT 2.605 2.530 2.835 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 4.910 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.505 0.300 2.735 0.765 ;
        RECT 0.000 -0.300 4.480 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.265 1.290 1.495 3.325 ;
        RECT 2.945 1.290 3.175 1.985 ;
        RECT 0.245 1.055 3.175 1.290 ;
        RECT 0.245 0.805 0.475 1.055 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and2_1
MACRO gf180mcu_fd_sc_mcu7t5v0__and2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.040 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.024000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.660 1.065 1.020 2.240 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.024000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.770 1.515 2.130 3.370 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.071900 ;
    PORT
      LAYER Metal1 ;
        RECT 3.420 0.550 3.830 3.355 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.040 4.220 ;
        RECT 0.260 2.545 0.490 3.620 ;
        RECT 2.520 2.530 2.750 3.620 ;
        RECT 4.560 2.530 4.790 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 5.470 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 5.470 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.300 0.300 2.530 0.690 ;
        RECT 4.560 0.300 4.790 0.765 ;
        RECT 0.000 -0.300 5.040 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.280 1.165 1.510 3.355 ;
        RECT 2.960 1.165 3.190 1.755 ;
        RECT 1.280 0.930 3.190 1.165 ;
        RECT 1.280 0.780 1.510 0.930 ;
        RECT 0.195 0.550 1.510 0.780 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and2_2
MACRO gf180mcu_fd_sc_mcu7t5v0__and2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.055000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.030 1.210 3.515 1.560 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.055000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.540 1.800 4.125 2.150 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.069600 ;
    PORT
      LAYER Metal1 ;
        RECT 5.470 2.710 5.810 3.380 ;
        RECT 7.510 2.710 7.930 3.380 ;
        RECT 5.470 2.330 7.930 2.710 ;
        RECT 7.370 1.245 7.930 2.330 ;
        RECT 5.390 0.920 7.930 1.245 ;
        RECT 5.390 0.825 5.730 0.920 ;
        RECT 7.370 0.550 7.930 0.920 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 9.520 4.220 ;
        RECT 0.245 2.530 0.475 3.620 ;
        RECT 2.285 3.040 2.515 3.620 ;
        RECT 4.325 3.040 4.555 3.620 ;
        RECT 6.545 3.040 6.775 3.620 ;
        RECT 8.585 2.530 8.815 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 9.950 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 0.905 ;
        RECT 4.325 0.300 4.555 0.765 ;
        RECT 6.510 0.300 6.850 0.640 ;
        RECT 8.805 0.300 9.035 0.905 ;
        RECT 0.000 -0.300 9.520 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.210 2.760 1.550 3.380 ;
        RECT 3.250 2.760 3.590 3.380 ;
        RECT 1.210 2.530 4.995 2.760 ;
        RECT 4.765 1.815 4.995 2.530 ;
        RECT 4.765 1.585 7.005 1.815 ;
        RECT 4.765 1.230 4.995 1.585 ;
        RECT 3.865 0.995 4.995 1.230 ;
        RECT 3.865 0.825 4.095 0.995 ;
        RECT 2.265 0.595 4.095 0.825 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and2_4
MACRO gf180mcu_fd_sc_mcu7t5v0__and3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.495500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.540 1.770 1.570 2.150 ;
        RECT 1.250 1.120 1.570 1.770 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.495500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 1.120 2.120 2.415 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.495500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.360 1.120 2.910 2.415 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.875600 ;
    PORT
      LAYER Metal1 ;
        RECT 4.570 0.650 5.010 3.380 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.600 4.220 ;
        RECT 1.210 3.285 1.550 3.620 ;
        RECT 3.745 2.530 3.975 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 6.030 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.645 0.300 3.875 1.090 ;
        RECT 0.000 -0.300 5.600 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 3.055 0.530 3.340 ;
        RECT 2.230 3.055 2.570 3.340 ;
        RECT 0.190 2.825 3.415 3.055 ;
        RECT 3.185 1.800 3.415 2.825 ;
        RECT 3.185 1.460 4.315 1.800 ;
        RECT 0.190 0.805 0.530 1.035 ;
        RECT 3.185 0.805 3.415 1.460 ;
        RECT 0.190 0.575 3.415 0.805 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and3_1
MACRO gf180mcu_fd_sc_mcu7t5v0__and3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.160 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.981500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.660 1.160 1.020 2.290 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.981500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.780 1.160 2.140 2.290 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.981500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.865 1.160 3.260 2.290 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.055600 ;
    PORT
      LAYER Metal1 ;
        RECT 4.480 0.650 4.950 3.380 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 6.160 4.220 ;
        RECT 1.320 3.160 1.550 3.620 ;
        RECT 3.360 3.160 3.590 3.620 ;
        RECT 5.580 2.530 5.810 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 6.590 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.590 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.360 0.300 3.590 0.765 ;
        RECT 5.600 0.300 5.830 0.765 ;
        RECT 0.000 -0.300 6.160 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.910 0.585 3.355 ;
        RECT 0.245 2.655 4.250 2.910 ;
        RECT 1.285 0.865 1.515 2.655 ;
        RECT 4.020 1.445 4.250 2.655 ;
        RECT 0.235 0.635 1.515 0.865 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and3_2
MACRO gf180mcu_fd_sc_mcu7t5v0__and3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.200 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.132000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.165 1.240 5.025 1.560 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.132000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.790 1.800 5.380 2.125 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.132000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.220 2.355 6.110 2.585 ;
        RECT 1.220 2.125 1.560 2.355 ;
        RECT 0.465 1.800 1.560 2.125 ;
        RECT 1.220 1.025 1.560 1.800 ;
        RECT 5.695 1.620 6.110 2.355 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.059200 ;
    PORT
      LAYER Metal1 ;
        RECT 7.550 2.725 7.890 3.340 ;
        RECT 9.590 2.725 9.990 3.340 ;
        RECT 7.550 2.385 9.990 2.725 ;
        RECT 9.610 1.100 9.990 2.385 ;
        RECT 7.250 0.870 9.990 1.100 ;
        RECT 7.250 0.810 7.590 0.870 ;
        RECT 9.545 0.550 9.990 0.870 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 11.200 4.220 ;
        RECT 0.245 2.530 0.475 3.620 ;
        RECT 2.230 3.285 2.570 3.620 ;
        RECT 4.270 3.285 4.610 3.620 ;
        RECT 6.530 3.285 6.870 3.620 ;
        RECT 8.570 3.285 8.910 3.620 ;
        RECT 10.665 2.530 10.895 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 11.630 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 11.630 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.325 0.300 0.555 0.695 ;
        RECT 6.185 0.300 6.415 0.765 ;
        RECT 8.370 0.300 8.710 0.640 ;
        RECT 10.665 0.300 10.895 0.905 ;
        RECT 0.000 -0.300 11.200 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.210 2.825 6.855 3.055 ;
        RECT 6.625 1.840 6.855 2.825 ;
        RECT 6.625 1.500 9.260 1.840 ;
        RECT 6.625 1.285 6.855 1.500 ;
        RECT 5.500 1.055 6.855 1.285 ;
        RECT 5.500 0.760 5.755 1.055 ;
        RECT 3.250 0.530 5.755 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and3_4
MACRO gf180mcu_fd_sc_mcu7t5v0__and4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.160 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.660 2.190 1.000 3.000 ;
        RECT 0.660 1.770 1.560 2.190 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.790 1.540 2.130 2.410 ;
        RECT 1.015 1.210 2.130 1.540 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.360 1.570 2.700 2.410 ;
        RECT 2.360 1.210 3.430 1.570 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.215 1.800 4.780 2.120 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.895400 ;
    PORT
      LAYER Metal1 ;
        RECT 5.660 0.610 6.030 3.350 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 6.160 4.220 ;
        RECT 0.250 3.285 0.590 3.620 ;
        RECT 2.290 3.285 2.630 3.620 ;
        RECT 4.550 3.285 4.890 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 6.590 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.590 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 4.505 0.300 4.845 1.035 ;
        RECT 0.000 -0.300 6.160 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.270 3.055 1.610 3.390 ;
        RECT 3.310 3.055 3.650 3.390 ;
        RECT 1.270 2.825 5.385 3.055 ;
        RECT 5.155 1.505 5.385 2.825 ;
        RECT 3.770 1.265 5.385 1.505 ;
        RECT 0.305 0.760 0.535 1.090 ;
        RECT 3.770 0.760 4.000 1.265 ;
        RECT 0.305 0.530 4.000 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and4_1
MACRO gf180mcu_fd_sc_mcu7t5v0__and4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.919500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.120 1.770 1.000 2.150 ;
        RECT 0.630 1.030 1.000 1.770 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.919500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.230 1.770 2.120 2.150 ;
        RECT 1.750 1.030 2.120 1.770 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.919500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.350 1.770 3.240 2.150 ;
        RECT 2.870 1.030 3.240 1.770 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.919500 ;
    PORT
      LAYER Metal1 ;
        RECT 3.470 1.770 4.595 2.150 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.060800 ;
    PORT
      LAYER Metal1 ;
        RECT 5.495 0.805 6.070 3.235 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.280 4.220 ;
        RECT 0.300 3.160 0.530 3.620 ;
        RECT 2.285 3.280 2.625 3.620 ;
        RECT 4.325 3.285 4.665 3.620 ;
        RECT 6.600 2.650 6.830 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 7.710 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 4.325 0.300 4.665 0.635 ;
        RECT 6.620 0.300 6.850 0.765 ;
        RECT 0.000 -0.300 7.280 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.260 2.790 5.230 3.020 ;
        RECT 5.000 1.095 5.230 2.790 ;
        RECT 3.845 0.865 5.230 1.095 ;
        RECT 3.845 0.780 4.075 0.865 ;
        RECT 0.235 0.550 4.075 0.780 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and4_2
MACRO gf180mcu_fd_sc_mcu7t5v0__and4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.440 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.884000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.215 1.770 2.570 2.135 ;
        RECT 2.340 1.675 2.570 1.770 ;
        RECT 2.340 1.445 3.870 1.675 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.884000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.825 1.905 7.545 2.135 ;
        RECT 5.420 1.800 7.545 1.905 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.884000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.960 1.215 2.050 1.385 ;
        RECT 6.830 1.220 7.170 1.380 ;
        RECT 4.005 1.215 7.170 1.220 ;
        RECT 0.960 0.990 7.170 1.215 ;
        RECT 0.960 0.985 4.235 0.990 ;
        RECT 0.960 0.680 3.890 0.985 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.884000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.140 2.365 8.280 2.595 ;
        RECT 0.140 1.770 0.985 2.365 ;
        RECT 7.960 1.645 8.280 2.365 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.939600 ;
    PORT
      LAYER Metal1 ;
        RECT 9.540 2.725 9.905 3.195 ;
        RECT 11.580 2.725 11.945 3.195 ;
        RECT 9.540 2.380 12.230 2.725 ;
        RECT 11.850 1.100 12.230 2.380 ;
        RECT 9.485 0.870 12.230 1.100 ;
        RECT 9.485 0.530 9.825 0.870 ;
        RECT 11.725 0.530 12.230 0.870 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 13.440 4.220 ;
        RECT 0.260 3.005 0.490 3.620 ;
        RECT 2.245 3.285 2.585 3.620 ;
        RECT 4.285 3.285 4.625 3.620 ;
        RECT 6.325 3.285 6.665 3.620 ;
        RECT 8.365 3.285 8.705 3.620 ;
        RECT 10.585 3.215 10.925 3.620 ;
        RECT 12.680 2.690 12.910 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 13.870 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.870 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.260 0.300 0.490 0.765 ;
        RECT 8.420 0.300 8.650 0.695 ;
        RECT 10.605 0.300 10.945 0.640 ;
        RECT 12.900 0.300 13.130 0.905 ;
        RECT 0.000 -0.300 13.440 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.185 2.825 9.090 3.055 ;
        RECT 8.860 1.755 9.090 2.825 ;
        RECT 8.860 1.525 11.550 1.755 ;
        RECT 8.860 1.155 9.090 1.525 ;
        RECT 7.960 0.925 9.090 1.155 ;
        RECT 7.960 0.760 8.190 0.925 ;
        RECT 4.285 0.530 8.190 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and4_4
MACRO gf180mcu_fd_sc_mcu7t5v0__antenna
  CLASS core ANTENNACELL ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__antenna ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.120 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.140 0.810 0.475 2.710 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 1.120 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 1.550 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 1.550 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.300 1.120 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__antenna
MACRO gf180mcu_fd_sc_mcu7t5v0__aoi21_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi21_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.099500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.775 1.770 2.680 2.150 ;
        RECT 2.340 1.160 2.680 1.770 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.099500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.115 1.770 1.010 2.150 ;
        RECT 0.660 1.160 1.010 1.770 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.913500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.910 1.770 3.815 2.150 ;
        RECT 3.475 1.160 3.815 1.770 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.145600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.240 0.870 1.545 2.725 ;
        RECT 1.240 0.550 2.580 0.870 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 4.480 4.220 ;
        RECT 3.525 2.690 3.755 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 4.910 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 0.765 ;
        RECT 3.625 0.300 3.855 0.765 ;
        RECT 0.000 -0.300 4.480 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 3.160 2.570 3.390 ;
        RECT 0.190 2.495 0.530 3.160 ;
        RECT 2.230 2.495 2.570 3.160 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi21_1
MACRO gf180mcu_fd_sc_mcu7t5v0__aoi21_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi21_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.145000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 1.240 6.725 1.560 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.145000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.290 1.800 6.725 2.120 ;
        RECT 3.290 1.400 3.630 1.800 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.893000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.580 1.800 2.280 2.125 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.081900 ;
    PORT
      LAYER Metal1 ;
        RECT 2.650 2.360 5.955 2.700 ;
        RECT 2.650 1.100 2.970 2.360 ;
        RECT 0.970 0.870 3.325 1.100 ;
        RECT 0.970 0.560 2.245 0.870 ;
        RECT 3.095 0.805 3.325 0.870 ;
        RECT 3.095 0.575 4.975 0.805 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.280 4.220 ;
        RECT 1.330 3.040 1.560 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 7.710 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.310 0.300 0.540 0.765 ;
        RECT 2.495 0.300 2.835 0.640 ;
        RECT 6.650 0.300 6.880 0.765 ;
        RECT 0.000 -0.300 7.280 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.310 2.760 0.540 3.380 ;
        RECT 1.800 3.095 6.880 3.325 ;
        RECT 1.800 2.760 2.035 3.095 ;
        RECT 0.310 2.530 2.035 2.760 ;
        RECT 6.650 2.435 6.880 3.095 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi21_2
MACRO gf180mcu_fd_sc_mcu7t5v0__aoi21_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi21_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.440 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.368000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 1.800 6.420 2.120 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.368000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.835 1.805 8.350 2.120 ;
        RECT 6.835 1.570 7.065 1.805 ;
        RECT 0.600 1.325 7.065 1.570 ;
        RECT 0.600 1.210 3.465 1.325 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.624000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.295 1.790 12.790 2.150 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.879200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.410 2.380 8.870 2.765 ;
        RECT 8.580 1.560 8.870 2.380 ;
        RECT 8.580 1.475 12.075 1.560 ;
        RECT 7.765 1.245 12.075 1.475 ;
        RECT 7.765 1.095 7.995 1.245 ;
        RECT 3.870 0.865 7.995 1.095 ;
        RECT 3.870 0.825 4.100 0.865 ;
        RECT 2.370 0.595 4.100 0.825 ;
        RECT 9.605 0.655 9.835 1.245 ;
        RECT 11.845 0.655 12.075 1.245 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 13.440 4.220 ;
        RECT 9.850 3.040 10.190 3.620 ;
        RECT 11.890 3.040 12.230 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 13.870 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.870 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.465 0.300 0.695 0.690 ;
        RECT 4.330 0.300 4.670 0.635 ;
        RECT 8.250 0.300 8.590 0.980 ;
        RECT 10.670 0.300 11.010 1.015 ;
        RECT 12.965 0.300 13.195 1.215 ;
        RECT 0.000 -0.300 13.440 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.445 3.160 9.565 3.390 ;
        RECT 0.445 2.540 0.675 3.160 ;
        RECT 9.235 2.760 9.565 3.160 ;
        RECT 10.870 2.760 11.210 3.380 ;
        RECT 12.910 2.760 13.250 3.380 ;
        RECT 9.235 2.530 13.250 2.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi21_4
MACRO gf180mcu_fd_sc_mcu7t5v0__aoi22_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi22_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.040 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.096500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.920 0.550 3.240 2.150 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.096500 ;
    PORT
      LAYER Metal1 ;
        RECT 3.480 1.800 4.545 2.150 ;
        RECT 3.480 0.550 3.800 1.800 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.096500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 0.550 2.120 2.150 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.096500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.610 1.770 1.570 2.150 ;
        RECT 0.610 1.085 1.005 1.770 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.055600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.350 2.380 3.890 2.710 ;
        RECT 2.350 0.585 2.680 2.380 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.040 4.220 ;
        RECT 1.330 3.040 1.560 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 5.470 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 5.470 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.310 0.300 0.540 0.725 ;
        RECT 4.390 0.300 4.620 0.905 ;
        RECT 0.000 -0.300 5.040 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.255 2.760 0.595 3.380 ;
        RECT 1.820 3.145 4.675 3.380 ;
        RECT 1.820 2.760 2.050 3.145 ;
        RECT 0.255 2.530 2.050 2.760 ;
        RECT 4.335 2.530 4.675 3.145 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi22_1
MACRO gf180mcu_fd_sc_mcu7t5v0__aoi22_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi22_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.960 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.193000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.690 1.210 8.380 1.570 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.193000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.950 1.800 8.380 2.120 ;
        RECT 4.950 1.400 5.235 1.800 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.193000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.650 1.030 2.090 1.590 ;
        RECT 0.940 0.610 2.090 1.030 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.193000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.620 1.820 4.030 2.120 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.139725 ;
    PORT
      LAYER Metal1 ;
        RECT 4.345 2.360 7.670 2.780 ;
        RECT 4.345 1.150 4.720 2.360 ;
        RECT 2.320 1.100 4.720 1.150 ;
        RECT 2.320 0.870 5.155 1.100 ;
        RECT 2.320 0.715 2.555 0.870 ;
        RECT 4.925 0.640 6.650 0.870 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 8.960 4.220 ;
        RECT 1.265 3.160 1.495 3.620 ;
        RECT 3.305 3.160 3.535 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 9.390 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.390 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 0.905 ;
        RECT 4.270 0.300 4.610 0.640 ;
        RECT 8.405 0.300 8.635 0.905 ;
        RECT 0.000 -0.300 8.960 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 2.760 0.530 3.380 ;
        RECT 2.230 2.760 2.570 3.380 ;
        RECT 3.795 3.130 8.690 3.365 ;
        RECT 3.795 2.760 4.025 3.130 ;
        RECT 0.190 2.530 4.025 2.760 ;
        RECT 8.350 2.475 8.690 3.130 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi22_2
MACRO gf180mcu_fd_sc_mcu7t5v0__aoi22_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi22_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.180 1.800 14.730 2.120 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.445 1.710 10.520 2.140 ;
        RECT 10.160 1.560 10.520 1.710 ;
        RECT 10.160 1.240 14.010 1.560 ;
        RECT 13.780 0.760 14.010 1.240 ;
        RECT 16.820 0.760 17.050 2.235 ;
        RECT 13.780 0.530 17.050 0.760 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.640 1.800 7.240 2.130 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.620 1.560 1.020 2.225 ;
        RECT 0.620 1.325 8.120 1.560 ;
        RECT 0.620 1.230 3.375 1.325 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.389000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.985 2.670 16.670 2.910 ;
        RECT 8.985 1.095 9.215 2.670 ;
        RECT 3.765 1.000 9.215 1.095 ;
        RECT 3.765 0.865 11.180 1.000 ;
        RECT 15.050 0.990 15.580 2.670 ;
        RECT 3.765 0.800 3.995 0.865 ;
        RECT 2.225 0.570 3.995 0.800 ;
        RECT 6.365 0.570 6.595 0.865 ;
        RECT 8.985 0.530 11.180 0.865 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 17.920 4.220 ;
        RECT 1.210 3.010 1.550 3.620 ;
        RECT 3.250 3.010 3.590 3.620 ;
        RECT 5.290 3.010 5.630 3.620 ;
        RECT 7.330 3.010 7.670 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 18.350 4.350 ;
        RECT -0.430 1.760 14.595 1.885 ;
        RECT 15.855 1.760 18.350 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 14.595 1.760 15.855 1.885 ;
        RECT -0.430 -0.430 18.350 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 0.695 ;
        RECT 4.270 0.300 4.610 0.635 ;
        RECT 8.350 0.300 8.690 0.635 ;
        RECT 12.845 0.300 13.075 0.730 ;
        RECT 17.365 0.300 17.595 0.730 ;
        RECT 0.000 -0.300 17.920 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 2.715 0.530 3.390 ;
        RECT 2.230 2.715 2.570 3.390 ;
        RECT 4.270 2.715 4.610 3.390 ;
        RECT 6.310 2.715 6.650 3.390 ;
        RECT 8.350 3.160 17.650 3.390 ;
        RECT 8.350 2.715 8.690 3.160 ;
        RECT 0.190 2.485 8.690 2.715 ;
        RECT 17.310 2.485 17.650 3.160 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi22_4
MACRO gf180mcu_fd_sc_mcu7t5v0__aoi211_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi211_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.033500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.770 1.770 2.690 2.150 ;
        RECT 1.770 1.230 2.150 1.770 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.033500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 1.160 1.000 2.190 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.886500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.920 2.850 4.010 3.310 ;
        RECT 2.920 1.730 3.220 2.850 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.886500 ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 1.770 4.950 2.150 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.259900 ;
    PORT
      LAYER Metal1 ;
        RECT 1.240 1.000 1.540 2.725 ;
        RECT 3.050 1.045 4.860 1.275 ;
        RECT 3.050 1.000 3.280 1.045 ;
        RECT 1.240 0.560 3.280 1.000 ;
        RECT 4.630 0.565 4.860 1.045 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.600 4.220 ;
        RECT 4.530 2.530 4.760 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 6.030 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 0.300 0.480 0.870 ;
        RECT 3.510 0.300 3.740 0.815 ;
        RECT 0.000 -0.300 5.600 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.250 3.150 2.520 3.380 ;
        RECT 0.250 2.530 0.480 3.150 ;
        RECT 2.290 2.530 2.520 3.150 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi211_1
MACRO gf180mcu_fd_sc_mcu7t5v0__aoi211_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi211_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.076000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.160 1.240 3.310 1.560 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.076000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.420 1.800 3.770 2.120 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.758000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.600 2.595 5.665 2.710 ;
        RECT 4.600 2.360 8.430 2.595 ;
        RECT 4.600 1.800 5.220 2.360 ;
        RECT 7.885 2.120 8.430 2.360 ;
        RECT 7.885 1.800 9.025 2.120 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.758000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.650 1.800 7.395 2.120 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.126800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.170 2.360 4.360 2.780 ;
        RECT 4.040 1.560 4.360 2.360 ;
        RECT 3.655 1.240 5.145 1.560 ;
        RECT 3.655 1.000 3.915 1.240 ;
        RECT 2.150 0.680 3.915 1.000 ;
        RECT 4.915 1.100 5.145 1.240 ;
        RECT 4.915 0.870 7.990 1.100 ;
        RECT 5.410 0.560 5.750 0.870 ;
        RECT 7.650 0.560 7.990 0.870 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 9.520 4.220 ;
        RECT 6.450 3.285 6.790 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 9.950 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 0.910 ;
        RECT 4.165 0.300 4.395 0.690 ;
        RECT 6.530 0.300 6.870 0.640 ;
        RECT 8.825 0.300 9.055 0.695 ;
        RECT 0.000 -0.300 9.520 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 3.160 6.140 3.390 ;
        RECT 0.245 2.500 0.475 3.160 ;
        RECT 5.910 3.055 6.140 3.160 ;
        RECT 8.725 3.055 8.955 3.390 ;
        RECT 5.910 2.825 8.955 3.055 ;
        RECT 8.725 2.500 8.955 2.825 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi211_2
MACRO gf180mcu_fd_sc_mcu7t5v0__aoi211_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi211_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.160 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.288000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.710 1.340 7.935 1.570 ;
        RECT 1.710 1.210 3.830 1.340 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.288000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.440 1.800 9.035 2.120 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.544000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.340 2.360 18.800 2.595 ;
        RECT 10.340 2.120 10.570 2.360 ;
        RECT 9.550 1.800 10.570 2.120 ;
        RECT 13.530 1.965 13.870 2.360 ;
        RECT 15.205 1.965 15.545 2.360 ;
        RECT 18.570 2.120 18.800 2.360 ;
        RECT 18.570 1.800 19.590 2.120 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.544000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.080 1.735 18.250 2.130 ;
        RECT 10.840 1.505 18.250 1.735 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.295200 ;
    PORT
      LAYER Metal1 ;
        RECT 0.980 2.360 8.340 2.680 ;
        RECT 0.980 1.185 1.210 2.360 ;
        RECT 0.980 0.955 1.420 1.185 ;
        RECT 8.505 1.100 18.740 1.275 ;
        RECT 1.190 0.930 1.420 0.955 ;
        RECT 4.480 1.045 18.740 1.100 ;
        RECT 4.480 0.930 8.735 1.045 ;
        RECT 1.190 0.870 8.735 0.930 ;
        RECT 1.190 0.700 4.710 0.870 ;
        RECT 2.900 0.530 3.240 0.700 ;
        RECT 6.980 0.575 7.320 0.870 ;
        RECT 10.360 0.775 10.700 1.045 ;
        RECT 13.040 0.775 13.380 1.045 ;
        RECT 15.720 0.775 16.060 1.045 ;
        RECT 18.400 0.775 18.740 1.045 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 20.160 4.220 ;
        RECT 11.700 3.285 12.040 3.620 ;
        RECT 16.975 3.285 17.315 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 20.590 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 20.590 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.620 0.300 0.960 0.710 ;
        RECT 4.940 0.300 5.280 0.640 ;
        RECT 9.020 0.300 9.360 0.765 ;
        RECT 11.700 0.300 12.040 0.710 ;
        RECT 14.380 0.300 14.720 0.765 ;
        RECT 17.060 0.300 17.400 0.765 ;
        RECT 19.575 0.300 19.805 1.060 ;
        RECT 0.000 -0.300 20.160 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.860 3.160 9.410 3.390 ;
        RECT 9.070 3.055 9.410 3.160 ;
        RECT 19.525 3.055 19.755 3.380 ;
        RECT 9.070 2.825 19.755 3.055 ;
        RECT 9.070 2.530 9.410 2.825 ;
        RECT 19.525 2.530 19.755 2.825 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi211_4
MACRO gf180mcu_fd_sc_mcu7t5v0__aoi221_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi221_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.160 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.033500 ;
    PORT
      LAYER Metal1 ;
        RECT 5.150 1.160 5.510 2.300 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.033500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.005 1.585 4.370 2.835 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.033500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.750 1.780 2.690 2.150 ;
        RECT 1.750 1.210 2.150 1.780 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.033500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.120 1.770 1.070 2.150 ;
        RECT 0.680 1.160 1.070 1.770 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.886500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.920 1.550 3.240 3.320 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.489200 ;
    PORT
      LAYER Metal1 ;
        RECT 4.600 1.205 4.920 2.865 ;
        RECT 2.950 0.975 4.920 1.205 ;
        RECT 2.950 0.905 3.180 0.975 ;
        RECT 2.150 0.675 3.180 0.905 ;
        RECT 4.600 0.905 4.920 0.975 ;
        RECT 4.600 0.675 5.980 0.905 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 6.160 4.220 ;
        RECT 1.365 3.160 1.595 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 6.590 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.590 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 0.815 ;
        RECT 3.670 0.300 4.010 0.745 ;
        RECT 0.000 -0.300 6.160 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.280 2.930 0.630 3.380 ;
        RECT 2.330 2.930 2.670 3.380 ;
        RECT 0.280 2.590 2.670 2.930 ;
        RECT 3.545 3.150 5.915 3.380 ;
        RECT 3.545 2.530 3.775 3.150 ;
        RECT 5.685 2.530 5.915 3.150 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi221_1
MACRO gf180mcu_fd_sc_mcu7t5v0__aoi221_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi221_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.880 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.978000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.080 1.790 12.050 2.120 ;
        RECT 9.080 1.550 9.310 1.790 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.978000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.570 1.225 12.050 1.560 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.978000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.125 1.910 7.815 2.140 ;
        RECT 5.650 1.800 7.815 1.910 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.978000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.525 1.785 3.270 2.150 ;
        RECT 3.040 1.680 3.270 1.785 ;
        RECT 3.040 1.450 5.390 1.680 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.870 1.325 2.810 1.555 ;
        RECT 2.580 1.220 2.810 1.325 ;
        RECT 5.770 1.220 8.310 1.560 ;
        RECT 2.580 1.210 8.310 1.220 ;
        RECT 2.580 0.990 6.000 1.210 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.496525 ;
    PORT
      LAYER Metal1 ;
        RECT 8.565 2.360 12.550 2.795 ;
        RECT 0.245 0.865 2.350 1.095 ;
        RECT 8.565 0.935 8.845 2.360 ;
        RECT 0.245 0.705 0.475 0.865 ;
        RECT 2.120 0.760 2.350 0.865 ;
        RECT 6.265 0.760 8.845 0.935 ;
        RECT 2.120 0.705 8.845 0.760 ;
        RECT 2.120 0.530 6.495 0.705 ;
        RECT 7.350 0.565 8.845 0.705 ;
        RECT 12.320 0.700 12.550 2.360 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 12.880 4.220 ;
        RECT 2.550 3.445 2.890 3.620 ;
        RECT 5.050 3.445 5.390 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 13.310 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.310 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.530 0.300 1.870 0.635 ;
        RECT 6.725 0.300 7.065 0.475 ;
        RECT 10.305 0.300 10.645 0.635 ;
        RECT 0.000 -0.300 12.880 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 3.215 2.290 3.350 ;
        RECT 5.855 3.215 12.505 3.365 ;
        RECT 0.345 3.135 12.505 3.215 ;
        RECT 0.345 3.120 6.195 3.135 ;
        RECT 0.345 2.460 0.575 3.120 ;
        RECT 2.075 2.985 6.195 3.120 ;
        RECT 1.310 2.525 7.410 2.755 ;
        RECT 8.105 2.460 8.335 3.135 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi221_2
MACRO gf180mcu_fd_sc_mcu7t5v0__aoi221_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi221_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.400 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.278000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.120 1.675 14.550 2.245 ;
        RECT 14.120 1.570 17.390 1.675 ;
        RECT 14.120 1.335 21.865 1.570 ;
        RECT 20.720 1.220 21.865 1.335 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.278000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.980 1.910 21.865 2.140 ;
        RECT 18.010 1.800 21.865 1.910 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.918000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.380 1.560 8.310 1.790 ;
        RECT 0.620 1.555 8.310 1.560 ;
        RECT 0.620 1.330 5.630 1.555 ;
        RECT 0.620 1.200 1.590 1.330 ;
        RECT 3.380 1.240 5.630 1.330 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.918000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.710 2.120 7.290 2.270 ;
        RECT 0.465 2.040 7.290 2.120 ;
        RECT 0.465 1.800 3.125 2.040 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.582000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.820 1.800 13.160 2.120 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.305500 ;
    PORT
      LAYER Metal1 ;
        RECT 13.530 2.680 21.050 2.910 ;
        RECT 13.530 1.560 13.880 2.680 ;
        RECT 8.905 1.325 13.880 1.560 ;
        RECT 5.880 1.105 13.880 1.325 ;
        RECT 1.820 0.960 3.080 1.100 ;
        RECT 0.190 0.870 3.080 0.960 ;
        RECT 0.190 0.730 2.050 0.870 ;
        RECT 2.850 0.780 3.080 0.870 ;
        RECT 5.880 1.095 16.470 1.105 ;
        RECT 5.880 0.780 6.110 1.095 ;
        RECT 2.850 0.545 6.110 0.780 ;
        RECT 8.555 0.765 8.785 1.095 ;
        RECT 11.110 0.530 11.450 1.095 ;
        RECT 13.530 0.875 16.470 1.095 ;
        RECT 13.530 0.530 13.870 0.875 ;
        RECT 16.240 0.780 16.470 0.875 ;
        RECT 18.460 0.870 20.470 1.105 ;
        RECT 18.460 0.780 18.690 0.870 ;
        RECT 16.240 0.545 18.690 0.780 ;
        RECT 20.240 0.775 20.470 0.870 ;
        RECT 20.240 0.545 22.040 0.775 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 22.400 4.220 ;
        RECT 0.240 2.530 0.580 3.620 ;
        RECT 2.335 3.040 2.565 3.620 ;
        RECT 4.375 3.040 4.605 3.620 ;
        RECT 6.415 3.040 6.645 3.620 ;
        RECT 8.455 3.040 8.685 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 22.830 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 22.830 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.280 0.300 2.620 0.640 ;
        RECT 6.360 0.300 6.700 0.795 ;
        RECT 10.045 0.300 10.275 0.795 ;
        RECT 12.285 0.300 12.515 0.795 ;
        RECT 15.570 0.300 15.910 0.640 ;
        RECT 19.650 0.300 19.990 0.640 ;
        RECT 0.000 -0.300 22.400 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.260 2.760 1.600 3.380 ;
        RECT 3.300 2.760 3.640 3.380 ;
        RECT 5.340 2.760 5.680 3.380 ;
        RECT 7.380 2.760 7.720 3.380 ;
        RECT 9.110 3.160 21.975 3.390 ;
        RECT 1.260 2.530 12.560 2.760 ;
        RECT 21.745 2.500 21.975 3.160 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi221_4
MACRO gf180mcu_fd_sc_mcu7t5v0__aoi222_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi222_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.072000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.840 2.330 7.720 2.710 ;
        RECT 6.840 1.230 7.180 2.330 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.072000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.140 2.330 6.040 2.710 ;
        RECT 5.720 1.535 6.040 2.330 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.072000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.350 1.770 3.800 2.150 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.072000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.040 1.770 4.950 2.150 ;
        RECT 4.040 1.105 4.360 1.770 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.072000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 0.550 2.120 2.235 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.072000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.480 1.770 1.560 2.150 ;
        RECT 1.240 0.550 1.560 1.770 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.756500 ;
    PORT
      LAYER Metal1 ;
        RECT 6.280 1.095 6.600 2.770 ;
        RECT 4.665 1.000 6.600 1.095 ;
        RECT 4.665 0.865 7.635 1.000 ;
        RECT 4.665 0.780 4.895 0.865 ;
        RECT 2.510 0.550 4.895 0.780 ;
        RECT 5.880 0.670 7.635 0.865 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.840 4.220 ;
        RECT 0.345 2.530 0.685 3.620 ;
        RECT 2.440 3.040 2.670 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 8.270 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.480 0.300 0.710 0.905 ;
        RECT 5.145 0.300 5.485 0.635 ;
        RECT 0.000 -0.300 7.840 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 2.760 1.705 3.380 ;
        RECT 3.095 3.095 7.635 3.325 ;
        RECT 1.365 2.530 4.500 2.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi222_1
MACRO gf180mcu_fd_sc_mcu7t5v0__aoi222_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi222_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.000 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.180000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.700 1.960 12.960 2.195 ;
        RECT 12.440 0.550 12.960 1.960 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.180000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.870 1.210 12.005 1.630 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.180000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.370 1.555 8.710 2.150 ;
        RECT 5.605 1.325 8.710 1.555 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.180000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.570 1.785 6.825 2.195 ;
        RECT 4.570 1.770 5.460 1.785 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.180000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.655 1.965 4.155 2.195 ;
        RECT 2.225 1.800 4.155 1.965 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.180000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 1.570 1.790 1.590 ;
        RECT 0.650 1.340 3.485 1.570 ;
        RECT 0.650 1.210 1.790 1.340 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.168800 ;
    PORT
      LAYER Metal1 ;
        RECT 9.050 2.440 13.485 2.670 ;
        RECT 9.050 1.095 9.470 2.440 ;
        RECT 2.020 0.970 9.470 1.095 ;
        RECT 0.225 0.865 9.470 0.970 ;
        RECT 0.225 0.740 2.250 0.865 ;
        RECT 4.925 0.845 5.265 0.865 ;
        RECT 9.050 0.790 9.470 0.865 ;
        RECT 13.255 0.570 13.485 2.440 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 14.000 4.220 ;
        RECT 0.225 2.530 0.565 3.620 ;
        RECT 2.320 3.040 2.550 3.620 ;
        RECT 4.360 3.040 4.590 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 14.430 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.430 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.455 0.300 2.795 0.635 ;
        RECT 7.065 0.300 7.405 0.635 ;
        RECT 11.160 0.300 11.500 0.635 ;
        RECT 0.000 -0.300 14.000 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.245 2.760 1.585 3.380 ;
        RECT 3.285 2.760 3.625 3.380 ;
        RECT 5.020 3.160 13.550 3.390 ;
        RECT 1.245 2.530 8.425 2.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi222_2
MACRO gf180mcu_fd_sc_mcu7t5v0__aoi222_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi222_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.320 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.408000 ;
    PORT
      LAYER Metal1 ;
        RECT 17.780 1.965 25.670 2.195 ;
        RECT 23.610 1.770 25.670 1.965 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.408000 ;
    PORT
      LAYER Metal1 ;
        RECT 17.535 1.325 23.110 1.615 ;
        RECT 17.535 1.160 18.430 1.325 ;
        RECT 20.405 1.220 22.490 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.408000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.945 1.565 10.160 2.150 ;
        RECT 16.605 1.565 16.835 2.025 ;
        RECT 8.945 1.335 16.835 1.565 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.408000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.415 1.800 16.255 2.120 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.408000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.320 1.760 8.515 2.150 ;
        RECT 7.320 1.565 7.620 1.760 ;
        RECT 0.710 1.335 7.620 1.565 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.408000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.585 1.800 7.090 2.120 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.940600 ;
    PORT
      LAYER Metal1 ;
        RECT 17.075 2.605 24.710 2.835 ;
        RECT 5.630 1.095 7.035 1.100 ;
        RECT 0.190 0.870 16.040 1.095 ;
        RECT 0.190 0.865 5.860 0.870 ;
        RECT 6.805 0.865 16.040 0.870 ;
        RECT 15.810 0.800 16.040 0.865 ;
        RECT 17.075 0.800 17.305 2.605 ;
        RECT 18.810 0.865 20.105 1.095 ;
        RECT 18.810 0.800 19.040 0.865 ;
        RECT 15.810 0.570 19.040 0.800 ;
        RECT 19.875 0.760 20.105 0.865 ;
        RECT 22.835 0.865 25.730 1.095 ;
        RECT 22.835 0.760 23.065 0.865 ;
        RECT 19.875 0.530 23.065 0.760 ;
        RECT 24.730 0.650 25.730 0.865 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 26.320 4.220 ;
        RECT 0.190 2.555 0.530 3.620 ;
        RECT 2.230 3.040 2.575 3.620 ;
        RECT 4.270 3.040 4.610 3.620 ;
        RECT 6.310 3.040 6.650 3.620 ;
        RECT 8.350 3.040 8.690 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 26.750 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 26.750 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.230 0.300 2.570 0.635 ;
        RECT 6.310 0.300 6.650 0.640 ;
        RECT 11.110 0.300 11.450 0.635 ;
        RECT 15.190 0.300 15.530 0.635 ;
        RECT 19.270 0.300 19.610 0.635 ;
        RECT 23.350 0.300 23.690 0.635 ;
        RECT 0.000 -0.300 26.320 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.210 2.760 1.550 3.380 ;
        RECT 3.250 2.760 3.590 3.380 ;
        RECT 5.290 2.760 5.630 3.380 ;
        RECT 7.330 2.760 7.670 3.380 ;
        RECT 9.070 3.160 25.730 3.390 ;
        RECT 1.210 2.530 16.550 2.760 ;
        RECT 25.390 2.555 25.730 3.160 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi222_4
MACRO gf180mcu_fd_sc_mcu7t5v0__buf_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 1.630 1.590 2.190 ;
        RECT 0.705 0.650 1.220 1.630 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.485 1.600 2.955 3.380 ;
        RECT 2.330 0.575 2.955 1.600 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 3.360 4.220 ;
        RECT 1.530 3.130 1.870 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 3.790 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 3.790 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.585 0.300 1.815 0.865 ;
        RECT 0.000 -0.300 3.360 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.815 0.630 3.390 ;
        RECT 0.245 2.580 2.255 2.815 ;
        RECT 0.245 0.800 0.475 2.580 ;
        RECT 1.970 1.830 2.255 2.580 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_1
MACRO gf180mcu_fd_sc_mcu7t5v0__buf_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 1.625 1.650 2.150 ;
        RECT 0.705 0.610 1.015 1.625 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal1 ;
        RECT 2.675 2.700 2.905 3.390 ;
        RECT 2.675 2.210 3.800 2.700 ;
        RECT 3.480 1.300 3.800 2.210 ;
        RECT 2.675 1.065 3.800 1.300 ;
        RECT 2.675 0.570 2.905 1.065 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 4.480 4.220 ;
        RECT 1.405 3.010 1.745 3.620 ;
        RECT 3.640 3.010 3.980 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 4.910 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.405 0.300 1.745 0.765 ;
        RECT 3.740 0.300 4.080 0.765 ;
        RECT 0.000 -0.300 4.480 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.625 0.475 3.390 ;
        RECT 0.245 2.390 2.130 2.625 ;
        RECT 0.245 0.570 0.475 2.390 ;
        RECT 1.900 1.890 2.130 2.390 ;
        RECT 1.900 1.550 3.240 1.890 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_2
MACRO gf180mcu_fd_sc_mcu7t5v0__buf_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 1.625 1.650 2.150 ;
        RECT 0.705 0.610 1.015 1.625 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal1 ;
        RECT 2.675 2.660 2.905 3.390 ;
        RECT 4.580 2.660 5.160 3.390 ;
        RECT 2.675 2.210 5.160 2.660 ;
        RECT 4.580 1.300 5.160 2.210 ;
        RECT 2.675 1.065 5.160 1.300 ;
        RECT 2.675 0.570 2.905 1.065 ;
        RECT 4.580 0.570 5.160 1.065 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.600 4.220 ;
        RECT 1.210 2.910 1.550 3.620 ;
        RECT 3.640 2.910 3.980 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 6.030 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.500 0.300 1.840 0.765 ;
        RECT 3.740 0.300 4.080 0.765 ;
        RECT 0.000 -0.300 5.600 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.625 0.475 3.390 ;
        RECT 0.245 2.390 2.130 2.625 ;
        RECT 0.245 0.570 0.475 2.390 ;
        RECT 1.900 1.890 2.130 2.390 ;
        RECT 1.900 1.550 4.175 1.890 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_3
MACRO gf180mcu_fd_sc_mcu7t5v0__buf_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.620 1.715 2.150 2.150 ;
        RECT 0.620 1.100 1.060 1.715 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal1 ;
        RECT 3.605 2.680 3.835 3.380 ;
        RECT 5.745 2.680 5.975 3.380 ;
        RECT 3.605 2.360 5.975 2.680 ;
        RECT 4.360 1.420 5.160 2.360 ;
        RECT 3.605 1.140 6.075 1.420 ;
        RECT 3.605 0.675 3.865 1.140 ;
        RECT 5.845 0.675 6.075 1.140 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.840 4.220 ;
        RECT 0.245 2.570 0.475 3.620 ;
        RECT 2.385 3.000 2.615 3.620 ;
        RECT 4.625 3.050 4.855 3.620 ;
        RECT 6.865 2.570 7.095 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 8.270 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 0.765 ;
        RECT 2.430 0.300 2.770 0.765 ;
        RECT 4.670 0.300 5.010 0.765 ;
        RECT 6.910 0.300 7.250 0.765 ;
        RECT 0.000 -0.300 7.840 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.265 2.760 1.495 3.380 ;
        RECT 1.265 2.530 2.905 2.760 ;
        RECT 2.670 2.025 2.905 2.530 ;
        RECT 2.670 1.685 4.095 2.025 ;
        RECT 5.585 1.685 6.810 2.025 ;
        RECT 2.670 1.250 2.905 1.685 ;
        RECT 1.365 1.015 2.905 1.250 ;
        RECT 1.365 0.675 1.595 1.015 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_4
MACRO gf180mcu_fd_sc_mcu7t5v0__buf_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.408000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 1.715 3.510 2.150 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal1 ;
        RECT 5.845 2.710 6.075 3.380 ;
        RECT 7.985 2.710 8.215 3.380 ;
        RECT 10.225 2.710 10.455 3.380 ;
        RECT 12.465 2.710 12.695 3.380 ;
        RECT 5.845 2.330 12.695 2.710 ;
        RECT 8.840 1.420 9.640 2.330 ;
        RECT 5.845 1.040 12.795 1.420 ;
        RECT 5.845 0.675 6.105 1.040 ;
        RECT 8.085 0.675 8.315 1.040 ;
        RECT 10.325 0.675 10.555 1.040 ;
        RECT 12.565 0.675 12.795 1.040 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 14.560 4.220 ;
        RECT 0.245 2.570 0.475 3.620 ;
        RECT 2.385 3.040 2.615 3.620 ;
        RECT 4.625 2.570 4.855 3.620 ;
        RECT 6.865 3.040 7.095 3.620 ;
        RECT 9.105 3.040 9.335 3.620 ;
        RECT 11.345 3.040 11.575 3.620 ;
        RECT 13.585 2.570 13.815 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 14.990 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 0.765 ;
        RECT 2.430 0.300 2.770 0.765 ;
        RECT 4.670 0.300 5.010 0.765 ;
        RECT 6.910 0.300 7.250 0.765 ;
        RECT 9.150 0.300 9.490 0.765 ;
        RECT 11.390 0.300 11.730 0.765 ;
        RECT 13.630 0.300 13.970 0.765 ;
        RECT 0.000 -0.300 14.560 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.265 2.760 1.495 3.380 ;
        RECT 3.505 2.760 3.735 3.380 ;
        RECT 1.265 2.530 4.315 2.760 ;
        RECT 3.980 2.025 4.315 2.530 ;
        RECT 3.980 1.685 8.270 2.025 ;
        RECT 10.340 1.685 13.540 2.030 ;
        RECT 3.980 1.250 4.315 1.685 ;
        RECT 1.365 1.015 4.315 1.250 ;
        RECT 1.365 0.675 1.595 1.015 ;
        RECT 3.605 0.675 3.835 1.015 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_8
MACRO gf180mcu_fd_sc_mcu7t5v0__buf_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.612000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.620 1.660 5.700 2.150 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal1 ;
        RECT 8.085 2.930 8.315 3.380 ;
        RECT 10.225 2.930 10.455 3.380 ;
        RECT 12.465 2.930 12.695 3.380 ;
        RECT 14.705 2.930 14.935 3.380 ;
        RECT 16.945 2.930 17.175 3.380 ;
        RECT 19.185 2.930 19.415 3.380 ;
        RECT 8.085 2.330 19.415 2.930 ;
        RECT 13.320 1.420 14.120 2.330 ;
        RECT 8.085 0.980 19.515 1.420 ;
        RECT 8.085 0.675 8.345 0.980 ;
        RECT 10.325 0.675 10.555 0.980 ;
        RECT 12.565 0.675 12.795 0.980 ;
        RECT 14.805 0.675 15.035 0.980 ;
        RECT 17.045 0.675 17.275 0.980 ;
        RECT 19.285 0.530 19.515 0.980 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 21.280 4.220 ;
        RECT 0.245 2.530 0.475 3.620 ;
        RECT 2.385 3.000 2.615 3.620 ;
        RECT 4.625 3.000 4.855 3.620 ;
        RECT 6.865 2.530 7.095 3.620 ;
        RECT 9.105 3.170 9.335 3.620 ;
        RECT 11.345 3.170 11.575 3.620 ;
        RECT 13.585 3.170 13.815 3.620 ;
        RECT 15.825 3.170 16.055 3.620 ;
        RECT 18.065 3.170 18.295 3.620 ;
        RECT 20.305 2.530 20.535 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 21.710 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.710 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 0.765 ;
        RECT 2.430 0.300 2.770 0.765 ;
        RECT 4.670 0.300 5.010 0.765 ;
        RECT 6.910 0.300 7.250 0.765 ;
        RECT 9.150 0.300 9.490 0.710 ;
        RECT 11.390 0.300 11.730 0.710 ;
        RECT 13.630 0.300 13.970 0.710 ;
        RECT 15.870 0.300 16.210 0.710 ;
        RECT 18.110 0.300 18.450 0.710 ;
        RECT 20.350 0.300 20.690 0.765 ;
        RECT 0.000 -0.300 21.280 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.265 2.760 1.495 3.380 ;
        RECT 3.505 2.760 3.735 3.380 ;
        RECT 5.745 2.760 5.975 3.380 ;
        RECT 1.265 2.530 6.495 2.760 ;
        RECT 6.260 2.025 6.495 2.530 ;
        RECT 6.260 1.685 12.805 2.025 ;
        RECT 14.625 1.685 20.260 2.030 ;
        RECT 6.260 1.250 6.495 1.685 ;
        RECT 1.365 1.015 6.495 1.250 ;
        RECT 1.365 0.675 1.595 1.015 ;
        RECT 3.605 0.675 3.835 1.015 ;
        RECT 5.845 0.675 6.075 1.015 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_12
MACRO gf180mcu_fd_sc_mcu7t5v0__buf_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.000 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 8.816000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.620 1.710 8.185 2.150 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.462399 ;
    PORT
      LAYER Metal1 ;
        RECT 10.325 2.810 10.555 3.380 ;
        RECT 12.465 2.810 12.695 3.380 ;
        RECT 14.705 2.810 14.935 3.380 ;
        RECT 16.945 2.810 17.175 3.380 ;
        RECT 19.185 2.810 19.415 3.380 ;
        RECT 21.425 2.810 21.655 3.380 ;
        RECT 23.665 2.810 23.895 3.380 ;
        RECT 25.905 2.810 26.135 3.380 ;
        RECT 10.325 2.230 26.135 2.810 ;
        RECT 17.750 1.510 18.650 2.230 ;
        RECT 10.325 0.930 26.235 1.510 ;
        RECT 10.325 0.675 10.585 0.930 ;
        RECT 12.565 0.675 12.795 0.930 ;
        RECT 14.805 0.675 15.035 0.930 ;
        RECT 17.045 0.675 17.275 0.930 ;
        RECT 19.285 0.675 19.515 0.930 ;
        RECT 21.525 0.675 21.755 0.930 ;
        RECT 23.765 0.675 23.995 0.930 ;
        RECT 26.005 0.675 26.235 0.930 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 28.000 4.220 ;
        RECT 0.245 2.530 0.475 3.620 ;
        RECT 2.385 3.000 2.615 3.620 ;
        RECT 4.625 3.000 4.855 3.620 ;
        RECT 6.865 3.000 7.095 3.620 ;
        RECT 9.105 2.530 9.335 3.620 ;
        RECT 11.345 3.040 11.575 3.620 ;
        RECT 13.585 3.040 13.815 3.620 ;
        RECT 15.825 3.040 16.055 3.620 ;
        RECT 18.065 3.040 18.295 3.620 ;
        RECT 20.305 3.040 20.535 3.620 ;
        RECT 22.545 3.040 22.775 3.620 ;
        RECT 24.785 3.040 25.015 3.620 ;
        RECT 27.025 2.530 27.255 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 28.430 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 28.430 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 0.765 ;
        RECT 2.430 0.300 2.770 0.765 ;
        RECT 4.670 0.300 5.010 0.765 ;
        RECT 6.910 0.300 7.250 0.765 ;
        RECT 9.150 0.300 9.490 0.765 ;
        RECT 11.390 0.300 11.730 0.700 ;
        RECT 13.630 0.300 13.970 0.700 ;
        RECT 15.870 0.300 16.210 0.700 ;
        RECT 18.110 0.300 18.450 0.700 ;
        RECT 20.350 0.300 20.690 0.700 ;
        RECT 22.590 0.300 22.930 0.700 ;
        RECT 24.830 0.300 25.170 0.700 ;
        RECT 27.070 0.300 27.410 0.765 ;
        RECT 0.000 -0.300 28.000 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.265 2.760 1.495 3.380 ;
        RECT 3.505 2.760 3.735 3.380 ;
        RECT 5.745 2.760 5.975 3.380 ;
        RECT 7.985 2.760 8.215 3.380 ;
        RECT 1.265 2.530 8.770 2.760 ;
        RECT 8.535 1.970 8.770 2.530 ;
        RECT 8.535 1.740 16.510 1.970 ;
        RECT 19.560 1.740 26.980 1.970 ;
        RECT 8.535 1.250 8.770 1.740 ;
        RECT 1.365 1.015 8.770 1.250 ;
        RECT 1.365 0.675 1.595 1.015 ;
        RECT 3.605 0.675 3.835 1.015 ;
        RECT 5.845 0.675 6.075 1.015 ;
        RECT 8.085 0.675 8.315 1.015 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_16
MACRO gf180mcu_fd_sc_mcu7t5v0__buf_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_20 ;
  ORIGIN 0.000 0.000 ;
  SIZE 34.720 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 11.020000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 1.740 9.900 2.150 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 11.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.565 3.000 12.795 3.380 ;
        RECT 14.705 3.000 14.935 3.380 ;
        RECT 16.945 3.000 17.175 3.380 ;
        RECT 19.185 3.000 19.415 3.380 ;
        RECT 21.425 3.000 21.655 3.380 ;
        RECT 23.665 3.000 23.895 3.380 ;
        RECT 25.905 3.000 26.135 3.380 ;
        RECT 28.145 3.000 28.375 3.380 ;
        RECT 30.385 3.000 30.615 3.380 ;
        RECT 32.625 3.000 32.855 3.380 ;
        RECT 12.565 2.270 32.855 3.000 ;
        RECT 22.230 1.510 23.130 2.270 ;
        RECT 12.565 0.865 32.955 1.510 ;
        RECT 12.565 0.675 12.825 0.865 ;
        RECT 14.805 0.675 15.035 0.865 ;
        RECT 17.045 0.675 17.275 0.865 ;
        RECT 19.285 0.675 19.515 0.865 ;
        RECT 21.525 0.675 21.755 0.865 ;
        RECT 23.765 0.675 23.995 0.865 ;
        RECT 26.005 0.675 26.235 0.865 ;
        RECT 28.245 0.675 28.475 0.865 ;
        RECT 30.485 0.675 30.715 0.865 ;
        RECT 32.725 0.675 32.955 0.865 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 34.720 4.220 ;
        RECT 0.245 2.530 0.475 3.620 ;
        RECT 2.385 3.000 2.615 3.620 ;
        RECT 4.625 3.000 4.855 3.620 ;
        RECT 6.865 3.000 7.095 3.620 ;
        RECT 9.105 3.000 9.335 3.620 ;
        RECT 11.345 2.530 11.575 3.620 ;
        RECT 13.585 3.230 13.815 3.620 ;
        RECT 15.825 3.230 16.055 3.620 ;
        RECT 18.065 3.230 18.295 3.620 ;
        RECT 20.305 3.230 20.535 3.620 ;
        RECT 22.545 3.230 22.775 3.620 ;
        RECT 24.785 3.230 25.015 3.620 ;
        RECT 27.025 3.230 27.255 3.620 ;
        RECT 29.265 3.230 29.495 3.620 ;
        RECT 31.505 3.230 31.735 3.620 ;
        RECT 33.745 2.530 33.975 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 35.150 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 35.150 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.160 ;
        RECT 2.485 0.300 2.715 0.960 ;
        RECT 4.725 0.300 4.955 0.960 ;
        RECT 6.965 0.300 7.195 0.960 ;
        RECT 9.205 0.300 9.435 0.960 ;
        RECT 11.445 0.300 11.675 0.960 ;
        RECT 13.630 0.300 13.970 0.635 ;
        RECT 15.870 0.300 16.210 0.635 ;
        RECT 18.110 0.300 18.450 0.635 ;
        RECT 20.350 0.300 20.690 0.635 ;
        RECT 22.590 0.300 22.930 0.635 ;
        RECT 24.830 0.300 25.170 0.635 ;
        RECT 27.070 0.300 27.410 0.635 ;
        RECT 29.310 0.300 29.650 0.635 ;
        RECT 31.550 0.300 31.890 0.635 ;
        RECT 33.845 0.300 34.075 1.160 ;
        RECT 0.000 -0.300 34.720 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 2.760 1.595 3.380 ;
        RECT 3.505 2.760 3.735 3.380 ;
        RECT 5.745 2.760 5.975 3.380 ;
        RECT 7.985 2.760 8.215 3.380 ;
        RECT 10.225 2.760 10.680 3.380 ;
        RECT 1.365 2.530 10.680 2.760 ;
        RECT 10.225 1.970 10.680 2.530 ;
        RECT 10.225 1.740 21.570 1.970 ;
        RECT 23.680 1.740 33.600 1.970 ;
        RECT 10.225 1.420 10.680 1.740 ;
        RECT 1.365 1.190 10.680 1.420 ;
        RECT 1.365 0.675 1.595 1.190 ;
        RECT 3.605 0.675 3.835 1.190 ;
        RECT 5.845 0.675 6.075 1.190 ;
        RECT 8.085 0.675 8.315 1.190 ;
        RECT 10.325 0.675 10.680 1.190 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_20
MACRO gf180mcu_fd_sc_mcu7t5v0__bufz_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__bufz_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.052000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.870 2.360 2.190 2.680 ;
        RECT 1.780 1.650 2.190 2.360 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.526000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.600 1.795 6.330 2.120 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 6.770 2.920 7.710 3.380 ;
        RECT 7.180 1.000 7.710 2.920 ;
        RECT 6.770 0.600 7.710 1.000 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.840 4.220 ;
        RECT 1.365 3.065 1.595 3.620 ;
        RECT 6.005 3.015 6.235 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 8.270 4.350 ;
        RECT -0.430 1.760 3.175 1.885 ;
        RECT 4.595 1.760 8.270 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 3.175 1.760 4.595 1.885 ;
        RECT -0.430 -0.430 8.270 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.760 ;
        RECT 6.225 0.300 6.455 0.790 ;
        RECT 0.000 -0.300 7.840 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 1.240 0.575 3.370 ;
        RECT 2.290 3.160 5.235 3.390 ;
        RECT 2.630 2.480 3.175 2.740 ;
        RECT 2.630 1.240 2.860 2.480 ;
        RECT 3.650 2.170 3.910 2.930 ;
        RECT 0.190 1.005 2.860 1.240 ;
        RECT 3.090 1.880 3.910 2.170 ;
        RECT 0.190 0.530 0.530 1.005 ;
        RECT 3.090 0.760 3.320 1.880 ;
        RECT 4.140 1.220 4.370 3.160 ;
        RECT 4.920 2.590 5.235 3.160 ;
        RECT 4.920 2.360 6.855 2.590 ;
        RECT 6.625 1.880 6.855 2.360 ;
        RECT 3.760 0.990 4.370 1.220 ;
        RECT 4.885 1.335 6.950 1.565 ;
        RECT 4.885 0.760 5.115 1.335 ;
        RECT 2.340 0.530 5.115 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__bufz_1
MACRO gf180mcu_fd_sc_mcu7t5v0__bufz_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__bufz_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.400 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.929000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.545 1.780 1.630 2.265 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.079500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.920 1.815 6.085 2.235 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.037400 ;
    PORT
      LAYER Metal1 ;
        RECT 6.805 0.600 7.160 3.380 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 8.400 4.220 ;
        RECT 1.450 3.260 1.790 3.620 ;
        RECT 5.830 3.220 6.170 3.620 ;
        RECT 7.870 2.530 8.210 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 8.830 4.350 ;
        RECT -0.430 1.760 2.875 1.885 ;
        RECT 4.530 1.760 8.830 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 2.875 1.760 4.530 1.885 ;
        RECT -0.430 -0.430 8.830 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.640 ;
        RECT 5.685 0.300 5.915 0.900 ;
        RECT 7.925 0.300 8.155 0.900 ;
        RECT 0.000 -0.300 8.400 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.700 3.160 5.175 3.390 ;
        RECT 0.420 2.780 2.130 3.010 ;
        RECT 4.460 2.930 5.175 3.160 ;
        RECT 1.900 2.520 2.130 2.780 ;
        RECT 1.900 2.235 3.650 2.520 ;
        RECT 1.900 1.325 2.130 2.235 ;
        RECT 3.890 2.005 4.230 2.930 ;
        RECT 0.190 1.095 2.130 1.325 ;
        RECT 2.485 1.775 4.230 2.005 ;
        RECT 4.460 2.700 6.565 2.930 ;
        RECT 0.190 0.865 0.530 1.095 ;
        RECT 2.485 0.760 2.715 1.775 ;
        RECT 4.460 1.545 4.690 2.700 ;
        RECT 6.335 1.900 6.565 2.700 ;
        RECT 3.770 1.315 4.690 1.545 ;
        RECT 5.125 1.355 6.510 1.585 ;
        RECT 3.770 0.990 4.110 1.315 ;
        RECT 5.125 0.760 5.355 1.355 ;
        RECT 2.485 0.530 5.355 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__bufz_2
MACRO gf180mcu_fd_sc_mcu7t5v0__bufz_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__bufz_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.200 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.929000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.545 1.775 1.630 2.185 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.658000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.090 1.800 7.275 2.120 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.915200 ;
    PORT
      LAYER Metal1 ;
        RECT 8.460 2.770 8.800 3.390 ;
        RECT 10.500 2.770 10.840 3.390 ;
        RECT 8.460 2.540 11.070 2.770 ;
        RECT 10.740 1.135 11.070 2.540 ;
        RECT 8.340 0.865 11.070 1.135 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 11.200 4.220 ;
        RECT 1.450 3.260 1.790 3.620 ;
        RECT 5.220 3.285 5.560 3.620 ;
        RECT 7.260 3.285 7.600 3.620 ;
        RECT 9.480 3.285 9.820 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.035 11.630 4.350 ;
        RECT -0.430 1.760 2.875 2.035 ;
        RECT 4.715 1.760 11.630 2.035 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 2.875 1.760 4.715 2.035 ;
        RECT -0.430 -0.430 11.630 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.655 ;
        RECT 4.670 0.300 5.010 0.475 ;
        RECT 7.220 0.300 7.560 0.635 ;
        RECT 9.550 0.300 9.890 0.635 ;
        RECT 0.000 -0.300 11.200 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.870 3.160 4.825 3.390 ;
        RECT 0.420 2.780 2.155 3.010 ;
        RECT 1.925 2.520 2.155 2.780 ;
        RECT 1.925 2.235 3.650 2.520 ;
        RECT 1.925 1.325 2.155 2.235 ;
        RECT 3.890 2.005 4.230 2.930 ;
        RECT 0.190 1.095 2.155 1.325 ;
        RECT 2.485 1.775 4.230 2.005 ;
        RECT 4.595 2.805 4.825 3.160 ;
        RECT 6.240 2.805 6.580 3.390 ;
        RECT 4.595 2.575 7.855 2.805 ;
        RECT 0.190 0.850 0.530 1.095 ;
        RECT 2.485 0.760 2.715 1.775 ;
        RECT 4.595 1.545 4.825 2.575 ;
        RECT 7.625 2.195 7.855 2.575 ;
        RECT 7.625 1.965 10.370 2.195 ;
        RECT 3.770 1.315 4.825 1.545 ;
        RECT 7.785 1.365 10.490 1.595 ;
        RECT 3.770 1.140 4.110 1.315 ;
        RECT 7.785 1.095 8.015 1.365 ;
        RECT 5.920 0.935 8.015 1.095 ;
        RECT 4.215 0.865 8.015 0.935 ;
        RECT 4.215 0.760 6.370 0.865 ;
        RECT 2.485 0.705 6.370 0.760 ;
        RECT 2.485 0.530 4.440 0.705 ;
        RECT 5.920 0.585 6.370 0.705 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__bufz_3
MACRO gf180mcu_fd_sc_mcu7t5v0__bufz_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__bufz_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.320 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.929000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 1.770 1.590 2.150 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.159000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.130 1.770 7.190 2.150 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.074800 ;
    PORT
      LAYER Metal1 ;
        RECT 8.350 2.800 8.690 3.380 ;
        RECT 10.390 2.800 10.730 3.380 ;
        RECT 8.350 2.760 10.730 2.800 ;
        RECT 8.350 2.520 11.110 2.760 ;
        RECT 10.730 1.135 11.110 2.520 ;
        RECT 8.160 0.865 11.110 1.135 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 12.320 4.220 ;
        RECT 1.450 3.260 1.790 3.620 ;
        RECT 5.290 3.285 5.630 3.620 ;
        RECT 7.330 3.285 7.670 3.620 ;
        RECT 9.370 3.285 9.710 3.620 ;
        RECT 11.410 3.285 11.750 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.035 12.750 4.350 ;
        RECT -0.430 1.760 2.875 2.035 ;
        RECT 4.715 1.760 12.750 2.035 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 2.875 1.760 4.715 2.035 ;
        RECT -0.430 -0.430 12.750 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.655 ;
        RECT 4.670 0.300 5.010 0.475 ;
        RECT 7.130 0.300 7.470 0.635 ;
        RECT 9.370 0.300 9.710 0.635 ;
        RECT 11.610 0.300 11.950 0.635 ;
        RECT 0.000 -0.300 12.320 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.870 3.160 4.825 3.390 ;
        RECT 0.420 2.780 2.155 3.010 ;
        RECT 1.925 2.520 2.155 2.780 ;
        RECT 1.925 2.235 3.650 2.520 ;
        RECT 1.925 1.325 2.155 2.235 ;
        RECT 3.890 2.005 4.230 2.930 ;
        RECT 0.190 1.095 2.155 1.325 ;
        RECT 2.485 1.775 4.230 2.005 ;
        RECT 4.595 2.760 4.825 3.160 ;
        RECT 6.310 2.760 6.650 3.380 ;
        RECT 4.595 2.530 7.745 2.760 ;
        RECT 0.190 0.850 0.530 1.095 ;
        RECT 2.485 0.760 2.715 1.775 ;
        RECT 4.595 1.545 4.825 2.530 ;
        RECT 7.515 2.195 7.745 2.530 ;
        RECT 7.515 1.965 10.150 2.195 ;
        RECT 3.770 1.315 4.825 1.545 ;
        RECT 7.515 1.365 10.150 1.595 ;
        RECT 3.770 1.140 4.110 1.315 ;
        RECT 7.515 1.095 7.745 1.365 ;
        RECT 5.695 0.935 7.745 1.095 ;
        RECT 4.215 0.865 7.745 0.935 ;
        RECT 4.215 0.760 5.945 0.865 ;
        RECT 2.485 0.705 5.945 0.760 ;
        RECT 2.485 0.530 4.440 0.705 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__bufz_4
MACRO gf180mcu_fd_sc_mcu7t5v0__bufz_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__bufz_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.040 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.929000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.545 1.775 1.675 2.185 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.318000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.075 1.800 9.430 2.120 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.149600 ;
    PORT
      LAYER Metal1 ;
        RECT 10.390 2.765 10.730 3.380 ;
        RECT 12.430 2.765 12.770 3.380 ;
        RECT 14.470 2.765 14.810 3.380 ;
        RECT 16.510 2.765 16.850 3.380 ;
        RECT 10.390 2.425 16.850 2.765 ;
        RECT 13.420 1.135 14.070 2.425 ;
        RECT 10.400 0.865 17.550 1.135 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 19.040 4.220 ;
        RECT 1.450 3.260 1.790 3.620 ;
        RECT 5.290 3.285 5.630 3.620 ;
        RECT 7.330 3.285 7.670 3.620 ;
        RECT 9.370 3.285 9.710 3.620 ;
        RECT 11.410 3.285 11.750 3.620 ;
        RECT 13.450 3.285 13.790 3.620 ;
        RECT 15.490 3.285 15.830 3.620 ;
        RECT 17.530 3.285 17.870 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.035 19.470 4.350 ;
        RECT -0.430 1.760 2.875 2.035 ;
        RECT 4.715 1.760 19.470 2.035 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 2.875 1.760 4.715 2.035 ;
        RECT -0.430 -0.430 19.470 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.655 ;
        RECT 4.670 0.300 5.010 0.475 ;
        RECT 7.130 0.300 7.470 0.635 ;
        RECT 9.370 0.300 9.710 0.635 ;
        RECT 11.610 0.300 11.950 0.635 ;
        RECT 13.850 0.300 14.190 0.635 ;
        RECT 16.090 0.300 16.430 0.635 ;
        RECT 18.330 0.300 18.670 0.635 ;
        RECT 0.000 -0.300 19.040 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.680 3.160 4.825 3.390 ;
        RECT 0.420 2.780 2.155 3.010 ;
        RECT 1.925 2.520 2.155 2.780 ;
        RECT 1.925 2.235 3.650 2.520 ;
        RECT 1.925 1.325 2.155 2.235 ;
        RECT 3.890 2.005 4.230 2.930 ;
        RECT 0.190 1.095 2.155 1.325 ;
        RECT 3.205 1.775 4.230 2.005 ;
        RECT 4.595 2.760 4.825 3.160 ;
        RECT 6.365 2.760 6.595 3.380 ;
        RECT 8.405 2.760 8.635 3.380 ;
        RECT 4.595 2.530 9.985 2.760 ;
        RECT 0.190 0.850 0.530 1.095 ;
        RECT 3.205 0.760 3.435 1.775 ;
        RECT 4.595 1.545 4.825 2.530 ;
        RECT 9.755 2.195 9.985 2.530 ;
        RECT 9.755 1.965 12.260 2.195 ;
        RECT 15.050 1.965 17.430 2.195 ;
        RECT 3.770 1.315 4.825 1.545 ;
        RECT 9.755 1.365 12.520 1.595 ;
        RECT 15.415 1.365 17.990 1.595 ;
        RECT 3.770 1.140 4.110 1.315 ;
        RECT 9.755 1.095 9.985 1.365 ;
        RECT 5.695 0.935 9.985 1.095 ;
        RECT 4.215 0.865 9.985 0.935 ;
        RECT 4.215 0.760 5.945 0.865 ;
        RECT 2.390 0.705 5.945 0.760 ;
        RECT 2.390 0.530 4.440 0.705 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__bufz_8
MACRO gf180mcu_fd_sc_mcu7t5v0__bufz_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__bufz_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.760 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.929000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.370 1.770 1.590 2.150 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.477000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.125 1.770 11.480 2.150 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.224400 ;
    PORT
      LAYER Metal1 ;
        RECT 12.630 2.970 12.970 3.380 ;
        RECT 14.670 2.970 15.010 3.380 ;
        RECT 16.710 2.970 17.050 3.380 ;
        RECT 18.750 2.970 19.090 3.380 ;
        RECT 20.790 2.970 21.130 3.380 ;
        RECT 22.830 2.970 23.170 3.380 ;
        RECT 12.630 2.530 23.170 2.970 ;
        RECT 17.900 1.135 18.500 2.530 ;
        RECT 12.730 0.865 24.270 1.135 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 25.760 4.220 ;
        RECT 1.450 3.260 1.790 3.620 ;
        RECT 5.490 3.040 5.830 3.620 ;
        RECT 7.530 3.040 7.870 3.620 ;
        RECT 9.570 3.040 9.910 3.620 ;
        RECT 11.610 3.040 11.950 3.620 ;
        RECT 13.650 3.285 13.990 3.620 ;
        RECT 15.690 3.285 16.030 3.620 ;
        RECT 17.730 3.285 18.070 3.620 ;
        RECT 19.770 3.285 20.110 3.620 ;
        RECT 21.810 3.285 22.150 3.620 ;
        RECT 23.850 3.040 24.190 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.035 26.190 4.350 ;
        RECT -0.430 1.760 2.875 2.035 ;
        RECT 4.715 1.760 26.190 2.035 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 2.875 1.760 4.715 2.035 ;
        RECT -0.430 -0.430 26.190 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.655 ;
        RECT 4.670 0.300 5.010 0.475 ;
        RECT 7.130 0.300 7.470 0.635 ;
        RECT 9.370 0.300 9.710 0.635 ;
        RECT 11.610 0.300 11.950 0.635 ;
        RECT 13.850 0.300 14.190 0.635 ;
        RECT 16.090 0.300 16.430 0.635 ;
        RECT 18.330 0.300 18.670 0.635 ;
        RECT 20.570 0.300 20.910 0.635 ;
        RECT 22.810 0.300 23.150 0.635 ;
        RECT 25.050 0.300 25.390 0.635 ;
        RECT 0.000 -0.300 25.760 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.685 3.160 4.825 3.390 ;
        RECT 0.420 2.780 2.135 3.010 ;
        RECT 1.905 2.520 2.135 2.780 ;
        RECT 1.905 2.235 3.650 2.520 ;
        RECT 1.905 1.325 2.135 2.235 ;
        RECT 3.890 2.005 4.230 2.930 ;
        RECT 0.190 1.095 2.135 1.325 ;
        RECT 2.485 1.775 4.230 2.005 ;
        RECT 4.595 2.760 4.825 3.160 ;
        RECT 6.510 2.760 6.850 3.380 ;
        RECT 8.550 2.760 8.890 3.380 ;
        RECT 10.590 2.760 10.930 3.380 ;
        RECT 4.595 2.530 12.010 2.760 ;
        RECT 0.190 0.850 0.530 1.095 ;
        RECT 2.485 0.760 2.715 1.775 ;
        RECT 4.595 1.545 4.825 2.530 ;
        RECT 11.780 2.195 12.010 2.530 ;
        RECT 11.780 1.965 17.490 2.195 ;
        RECT 19.330 1.965 23.705 2.195 ;
        RECT 3.770 1.315 4.825 1.545 ;
        RECT 11.780 1.365 16.875 1.595 ;
        RECT 19.010 1.365 23.705 1.595 ;
        RECT 3.770 1.140 4.110 1.315 ;
        RECT 11.780 1.095 12.010 1.365 ;
        RECT 5.695 0.935 12.010 1.095 ;
        RECT 4.215 0.865 12.010 0.935 ;
        RECT 4.215 0.760 5.945 0.865 ;
        RECT 2.485 0.705 5.945 0.760 ;
        RECT 2.485 0.530 4.440 0.705 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__bufz_12
MACRO gf180mcu_fd_sc_mcu7t5v0__bufz_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__bufz_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 32.480 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.898000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.370 1.770 1.590 2.150 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 8.548500 ;
    PORT
      LAYER Metal1 ;
        RECT 5.690 1.770 12.790 2.150 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 8.299200 ;
    PORT
      LAYER Metal1 ;
        RECT 14.950 3.055 15.290 3.380 ;
        RECT 16.990 3.055 17.330 3.380 ;
        RECT 19.030 3.055 19.370 3.380 ;
        RECT 21.070 3.055 21.410 3.380 ;
        RECT 23.130 3.055 23.450 3.380 ;
        RECT 25.150 3.055 25.490 3.380 ;
        RECT 27.190 3.055 27.530 3.380 ;
        RECT 29.230 3.055 29.570 3.380 ;
        RECT 14.950 2.505 29.570 3.055 ;
        RECT 22.230 1.095 23.130 2.505 ;
        RECT 14.970 0.865 30.990 1.095 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 32.480 4.220 ;
        RECT 1.450 3.260 1.790 3.620 ;
        RECT 5.290 3.040 5.630 3.620 ;
        RECT 7.330 3.040 7.670 3.620 ;
        RECT 9.370 3.040 9.710 3.620 ;
        RECT 11.710 3.040 12.050 3.620 ;
        RECT 13.930 2.530 14.270 3.620 ;
        RECT 15.970 3.285 16.310 3.620 ;
        RECT 18.010 3.285 18.350 3.620 ;
        RECT 20.050 3.285 20.390 3.620 ;
        RECT 22.090 3.285 22.430 3.620 ;
        RECT 24.130 3.285 24.470 3.620 ;
        RECT 26.170 3.285 26.510 3.620 ;
        RECT 28.210 3.285 28.550 3.620 ;
        RECT 30.305 2.530 30.535 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 2.035 32.910 4.350 ;
        RECT -0.430 1.760 2.875 2.035 ;
        RECT 4.745 1.760 32.910 2.035 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 2.875 1.760 4.745 2.035 ;
        RECT -0.430 -0.430 32.910 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.640 ;
        RECT 4.670 0.300 5.010 0.475 ;
        RECT 7.130 0.300 7.470 0.635 ;
        RECT 9.370 0.300 9.710 0.635 ;
        RECT 11.610 0.300 11.950 0.635 ;
        RECT 13.835 0.300 14.210 0.635 ;
        RECT 16.090 0.300 16.430 0.635 ;
        RECT 18.330 0.300 18.670 0.635 ;
        RECT 20.570 0.300 20.910 0.635 ;
        RECT 22.810 0.300 23.150 0.635 ;
        RECT 25.050 0.300 25.390 0.635 ;
        RECT 27.290 0.300 27.630 0.635 ;
        RECT 29.530 0.300 29.870 0.635 ;
        RECT 31.825 0.300 32.055 0.900 ;
        RECT 0.000 -0.300 32.480 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.730 3.160 5.060 3.390 ;
        RECT 0.420 2.780 2.125 3.010 ;
        RECT 1.895 2.520 2.125 2.780 ;
        RECT 1.895 2.235 3.650 2.520 ;
        RECT 1.895 1.325 2.125 2.235 ;
        RECT 3.890 2.005 4.230 2.930 ;
        RECT 0.190 1.095 2.125 1.325 ;
        RECT 2.485 1.775 4.230 2.005 ;
        RECT 4.830 2.760 5.060 3.160 ;
        RECT 6.310 2.760 6.650 3.380 ;
        RECT 8.350 2.760 8.690 3.380 ;
        RECT 10.545 2.760 10.885 3.380 ;
        RECT 12.790 2.760 13.130 3.380 ;
        RECT 4.830 2.530 13.615 2.760 ;
        RECT 0.190 0.865 0.530 1.095 ;
        RECT 2.485 0.760 2.715 1.775 ;
        RECT 4.830 1.545 5.060 2.530 ;
        RECT 13.270 2.230 13.615 2.530 ;
        RECT 13.270 2.000 21.920 2.230 ;
        RECT 23.630 2.000 30.080 2.230 ;
        RECT 3.770 1.315 5.060 1.545 ;
        RECT 13.350 1.360 21.450 1.590 ;
        RECT 23.490 1.360 31.520 1.590 ;
        RECT 3.770 1.140 4.110 1.315 ;
        RECT 13.350 1.095 13.640 1.360 ;
        RECT 6.010 0.935 13.640 1.095 ;
        RECT 4.215 0.865 13.640 0.935 ;
        RECT 4.215 0.760 6.350 0.865 ;
        RECT 2.485 0.705 6.350 0.760 ;
        RECT 2.485 0.530 4.440 0.705 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__bufz_16
MACRO gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.741000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 1.740 1.590 2.150 ;
        RECT 0.705 1.035 1.080 1.740 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.754600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.565 1.605 2.930 3.320 ;
        RECT 2.340 0.565 2.930 1.605 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 3.360 4.220 ;
        RECT 1.310 3.015 1.650 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 3.790 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 3.790 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.925 ;
        RECT 0.000 -0.300 3.360 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.755 0.575 3.380 ;
        RECT 0.245 2.520 2.270 2.755 ;
        RECT 0.245 0.565 0.475 2.520 ;
        RECT 1.930 1.880 2.270 2.520 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
MACRO gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.726000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 1.740 1.650 2.150 ;
        RECT 0.705 0.550 1.080 1.740 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.008600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.665 2.710 2.895 3.390 ;
        RECT 2.665 2.360 3.810 2.710 ;
        RECT 3.470 1.510 3.810 2.360 ;
        RECT 2.665 1.280 3.810 1.510 ;
        RECT 2.665 0.800 2.895 1.280 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 4.480 4.220 ;
        RECT 1.360 3.050 1.700 3.620 ;
        RECT 3.685 3.050 3.915 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 4.910 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.490 0.300 1.830 1.095 ;
        RECT 3.730 0.300 4.070 1.050 ;
        RECT 0.000 -0.300 4.480 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.820 0.475 3.390 ;
        RECT 0.245 2.590 2.215 2.820 ;
        RECT 0.245 0.805 0.475 2.590 ;
        RECT 1.890 2.040 2.215 2.590 ;
        RECT 1.890 1.740 3.210 2.040 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
MACRO gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.183000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.620 1.740 2.340 2.120 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.785 2.680 4.015 3.390 ;
        RECT 5.925 2.680 6.155 3.390 ;
        RECT 3.785 2.360 6.600 2.680 ;
        RECT 6.280 1.510 6.600 2.360 ;
        RECT 3.785 1.280 6.600 1.510 ;
        RECT 3.785 0.690 4.015 1.280 ;
        RECT 6.025 0.690 6.255 1.280 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.840 4.220 ;
        RECT 0.245 3.200 0.475 3.620 ;
        RECT 2.385 3.160 2.615 3.620 ;
        RECT 4.805 3.050 5.035 3.620 ;
        RECT 7.045 2.730 7.275 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 8.270 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 0.985 ;
        RECT 2.610 0.300 2.950 0.985 ;
        RECT 4.850 0.300 5.190 0.985 ;
        RECT 7.090 0.300 7.430 0.985 ;
        RECT 0.000 -0.300 7.840 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.265 2.820 1.495 3.390 ;
        RECT 1.265 2.590 3.185 2.820 ;
        RECT 2.955 2.040 3.185 2.590 ;
        RECT 2.955 1.740 5.945 2.040 ;
        RECT 2.955 1.500 3.185 1.740 ;
        RECT 1.365 1.270 3.185 1.500 ;
        RECT 1.365 0.690 1.595 1.270 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
MACRO gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.183000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.370 1.740 2.150 2.150 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.785 2.680 4.015 3.390 ;
        RECT 5.925 2.680 6.155 3.390 ;
        RECT 3.785 2.360 6.155 2.680 ;
        RECT 5.130 1.445 5.510 2.360 ;
        RECT 3.785 1.215 6.255 1.445 ;
        RECT 3.785 0.690 4.015 1.215 ;
        RECT 6.025 0.690 6.255 1.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.840 4.220 ;
        RECT 0.245 3.230 0.475 3.620 ;
        RECT 2.385 3.160 2.615 3.620 ;
        RECT 4.805 3.050 5.035 3.620 ;
        RECT 7.045 2.760 7.275 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 8.270 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 1.040 ;
        RECT 2.610 0.300 2.950 0.985 ;
        RECT 4.850 0.300 5.190 0.985 ;
        RECT 7.090 0.300 7.430 0.985 ;
        RECT 0.000 -0.300 7.840 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.265 2.760 1.495 3.380 ;
        RECT 1.265 2.530 3.175 2.760 ;
        RECT 2.945 2.025 3.175 2.530 ;
        RECT 2.945 1.685 4.830 2.025 ;
        RECT 5.765 1.685 6.935 2.025 ;
        RECT 2.945 1.500 3.175 1.685 ;
        RECT 1.365 1.270 3.175 1.500 ;
        RECT 1.365 0.740 1.595 1.270 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
MACRO gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.369000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 1.745 4.130 2.150 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.408000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.025 2.680 6.255 3.390 ;
        RECT 8.265 2.680 8.495 3.390 ;
        RECT 10.505 2.680 10.735 3.390 ;
        RECT 12.745 2.680 12.975 3.390 ;
        RECT 6.025 2.360 12.975 2.680 ;
        RECT 9.610 1.510 9.990 2.360 ;
        RECT 6.025 1.220 12.975 1.510 ;
        RECT 6.025 0.690 6.255 1.220 ;
        RECT 8.265 0.690 8.495 1.220 ;
        RECT 10.505 0.690 10.735 1.220 ;
        RECT 12.745 0.690 12.975 1.220 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 14.560 4.220 ;
        RECT 0.245 3.230 0.475 3.620 ;
        RECT 2.485 3.050 2.715 3.620 ;
        RECT 4.905 3.230 5.135 3.620 ;
        RECT 7.145 3.050 7.375 3.620 ;
        RECT 9.385 3.050 9.615 3.620 ;
        RECT 11.625 3.050 11.855 3.620 ;
        RECT 13.865 2.760 14.095 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 14.990 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 1.040 ;
        RECT 2.430 0.300 2.770 1.040 ;
        RECT 4.850 0.300 5.190 1.055 ;
        RECT 7.090 0.300 7.430 0.985 ;
        RECT 9.330 0.300 9.670 0.985 ;
        RECT 11.570 0.300 11.910 0.985 ;
        RECT 13.810 0.300 14.150 0.985 ;
        RECT 0.000 -0.300 14.560 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 2.760 1.595 3.390 ;
        RECT 3.605 2.760 3.835 3.390 ;
        RECT 1.365 2.530 4.655 2.760 ;
        RECT 4.425 1.975 4.655 2.530 ;
        RECT 4.425 1.740 8.920 1.975 ;
        RECT 10.530 1.740 13.720 2.040 ;
        RECT 4.425 1.500 4.655 1.740 ;
        RECT 1.365 1.270 4.655 1.500 ;
        RECT 1.365 0.740 1.595 1.270 ;
        RECT 3.605 0.740 3.835 1.270 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
MACRO gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.555000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.620 1.765 6.070 2.150 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.036000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.265 3.000 8.495 3.390 ;
        RECT 10.405 3.000 10.635 3.390 ;
        RECT 12.645 3.000 12.875 3.390 ;
        RECT 14.885 3.000 15.115 3.390 ;
        RECT 17.125 3.000 17.355 3.390 ;
        RECT 19.365 3.000 19.595 3.390 ;
        RECT 8.265 2.495 19.595 3.000 ;
        RECT 13.830 1.535 14.730 2.495 ;
        RECT 8.265 1.215 19.695 1.535 ;
        RECT 8.265 0.690 8.495 1.215 ;
        RECT 10.505 0.690 10.735 1.215 ;
        RECT 12.745 0.690 12.975 1.215 ;
        RECT 14.985 0.690 15.215 1.215 ;
        RECT 17.225 0.690 17.455 1.215 ;
        RECT 19.465 0.690 19.695 1.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 21.280 4.220 ;
        RECT 0.245 3.230 0.475 3.620 ;
        RECT 2.385 3.050 2.615 3.620 ;
        RECT 4.625 3.050 4.855 3.620 ;
        RECT 7.145 3.230 7.375 3.620 ;
        RECT 9.285 3.230 9.515 3.620 ;
        RECT 11.525 3.230 11.755 3.620 ;
        RECT 13.765 3.230 13.995 3.620 ;
        RECT 16.005 3.230 16.235 3.620 ;
        RECT 18.245 3.230 18.475 3.620 ;
        RECT 20.485 2.760 20.715 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 21.710 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.710 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 1.075 ;
        RECT 2.430 0.300 2.770 1.075 ;
        RECT 4.670 0.300 5.010 1.075 ;
        RECT 7.090 0.300 7.430 1.075 ;
        RECT 9.330 0.300 9.670 0.985 ;
        RECT 11.570 0.300 11.910 0.985 ;
        RECT 13.810 0.300 14.150 0.985 ;
        RECT 16.050 0.300 16.390 0.985 ;
        RECT 18.290 0.300 18.630 0.985 ;
        RECT 20.530 0.300 20.870 0.985 ;
        RECT 0.000 -0.300 21.280 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.265 2.760 1.495 3.390 ;
        RECT 3.505 2.760 3.735 3.390 ;
        RECT 5.745 2.760 5.975 3.390 ;
        RECT 1.265 2.530 6.595 2.760 ;
        RECT 6.365 2.065 6.595 2.530 ;
        RECT 6.365 1.765 13.090 2.065 ;
        RECT 15.390 1.765 20.430 2.065 ;
        RECT 6.365 1.535 6.595 1.765 ;
        RECT 1.310 1.305 6.595 1.535 ;
        RECT 1.310 0.845 1.650 1.305 ;
        RECT 3.550 0.845 3.890 1.305 ;
        RECT 5.790 0.845 6.130 1.305 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
MACRO gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.000 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.738000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.370 1.740 8.310 2.150 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 8.068800 ;
    PORT
      LAYER Metal1 ;
        RECT 10.505 3.000 10.735 3.390 ;
        RECT 12.645 3.000 12.875 3.390 ;
        RECT 14.885 3.000 15.115 3.390 ;
        RECT 17.125 3.000 17.355 3.390 ;
        RECT 19.365 3.000 19.595 3.390 ;
        RECT 21.605 3.000 21.835 3.390 ;
        RECT 23.845 3.000 24.075 3.390 ;
        RECT 26.085 3.000 26.315 3.390 ;
        RECT 10.505 2.420 26.315 3.000 ;
        RECT 17.985 1.535 18.885 2.420 ;
        RECT 10.505 1.215 26.415 1.535 ;
        RECT 10.505 0.690 10.735 1.215 ;
        RECT 12.745 0.690 12.975 1.215 ;
        RECT 14.985 0.690 15.215 1.215 ;
        RECT 17.225 0.690 17.455 1.215 ;
        RECT 19.465 0.690 19.695 1.215 ;
        RECT 21.705 0.690 21.935 1.215 ;
        RECT 23.945 0.690 24.175 1.215 ;
        RECT 26.185 0.690 26.415 1.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 28.000 4.220 ;
        RECT 0.245 3.230 0.475 3.620 ;
        RECT 2.385 3.050 2.615 3.620 ;
        RECT 4.625 3.050 4.855 3.620 ;
        RECT 6.865 3.050 7.095 3.620 ;
        RECT 9.385 3.190 9.615 3.620 ;
        RECT 11.525 3.230 11.755 3.620 ;
        RECT 13.765 3.230 13.995 3.620 ;
        RECT 16.005 3.230 16.235 3.620 ;
        RECT 18.245 3.230 18.475 3.620 ;
        RECT 20.485 3.230 20.715 3.620 ;
        RECT 22.725 3.230 22.955 3.620 ;
        RECT 24.965 3.230 25.195 3.620 ;
        RECT 27.205 2.760 27.435 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 28.430 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 28.430 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.430 0.300 2.770 1.040 ;
        RECT 4.670 0.300 5.010 1.040 ;
        RECT 6.910 0.300 7.250 1.040 ;
        RECT 9.330 0.300 9.670 0.960 ;
        RECT 11.570 0.300 11.910 0.985 ;
        RECT 13.810 0.300 14.150 0.985 ;
        RECT 16.050 0.300 16.390 0.985 ;
        RECT 18.290 0.300 18.630 0.985 ;
        RECT 20.530 0.300 20.870 0.985 ;
        RECT 22.770 0.300 23.110 0.985 ;
        RECT 25.010 0.300 25.350 0.985 ;
        RECT 27.250 0.300 27.590 0.985 ;
        RECT 0.000 -0.300 28.000 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.265 2.760 1.495 3.390 ;
        RECT 3.505 2.760 3.735 3.390 ;
        RECT 5.745 2.760 5.975 3.390 ;
        RECT 7.985 2.760 8.215 3.390 ;
        RECT 1.265 2.530 8.850 2.760 ;
        RECT 8.620 2.065 8.850 2.530 ;
        RECT 8.620 1.765 17.160 2.065 ;
        RECT 19.740 1.765 27.160 2.065 ;
        RECT 8.620 1.500 8.850 1.765 ;
        RECT 1.365 1.270 8.850 1.500 ;
        RECT 1.365 0.740 1.595 1.270 ;
        RECT 3.605 0.740 3.835 1.270 ;
        RECT 5.845 0.740 6.075 1.270 ;
        RECT 8.085 0.740 8.315 1.270 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
MACRO gf180mcu_fd_sc_mcu7t5v0__clkbuf_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 ;
  ORIGIN 0.000 0.000 ;
  SIZE 34.720 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.924000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 1.740 9.900 2.120 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 10.130000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.745 3.000 12.975 3.390 ;
        RECT 14.885 3.000 15.115 3.390 ;
        RECT 17.125 3.000 17.355 3.390 ;
        RECT 19.365 3.000 19.595 3.390 ;
        RECT 21.605 3.000 21.835 3.390 ;
        RECT 23.845 3.000 24.075 3.390 ;
        RECT 26.085 3.000 26.315 3.390 ;
        RECT 28.325 3.000 28.555 3.390 ;
        RECT 30.565 3.000 30.795 3.390 ;
        RECT 32.905 3.000 33.135 3.390 ;
        RECT 12.745 2.270 33.135 3.000 ;
        RECT 22.230 1.535 23.130 2.270 ;
        RECT 12.745 1.215 33.135 1.535 ;
        RECT 12.745 0.685 13.005 1.215 ;
        RECT 14.985 0.685 15.215 1.215 ;
        RECT 17.225 0.685 17.455 1.215 ;
        RECT 19.465 0.685 19.695 1.215 ;
        RECT 21.705 0.685 21.935 1.215 ;
        RECT 23.945 0.685 24.175 1.215 ;
        RECT 26.185 0.685 26.415 1.215 ;
        RECT 28.425 0.685 28.655 1.215 ;
        RECT 30.665 0.685 30.895 1.215 ;
        RECT 32.905 0.685 33.135 1.215 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 34.720 4.220 ;
        RECT 0.245 3.230 0.475 3.620 ;
        RECT 2.385 3.050 2.615 3.620 ;
        RECT 4.625 3.050 4.855 3.620 ;
        RECT 6.865 3.050 7.095 3.620 ;
        RECT 9.105 3.050 9.335 3.620 ;
        RECT 11.625 3.230 11.855 3.620 ;
        RECT 13.765 3.230 13.995 3.620 ;
        RECT 16.005 3.230 16.235 3.620 ;
        RECT 18.245 3.230 18.475 3.620 ;
        RECT 20.485 3.230 20.715 3.620 ;
        RECT 22.725 3.230 22.955 3.620 ;
        RECT 24.965 3.230 25.195 3.620 ;
        RECT 27.205 3.230 27.435 3.620 ;
        RECT 29.445 3.230 29.675 3.620 ;
        RECT 31.685 3.230 31.915 3.620 ;
        RECT 34.025 2.710 34.255 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 35.150 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 35.150 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.485 0.300 2.715 1.040 ;
        RECT 4.725 0.300 4.955 1.040 ;
        RECT 6.965 0.300 7.195 1.040 ;
        RECT 9.205 0.300 9.435 1.040 ;
        RECT 11.445 0.300 11.675 1.040 ;
        RECT 13.810 0.300 14.150 0.985 ;
        RECT 16.050 0.300 16.390 0.985 ;
        RECT 18.290 0.300 18.630 0.985 ;
        RECT 20.530 0.300 20.870 0.985 ;
        RECT 22.770 0.300 23.110 0.985 ;
        RECT 25.010 0.300 25.350 0.985 ;
        RECT 27.250 0.300 27.590 0.985 ;
        RECT 29.490 0.300 29.830 0.985 ;
        RECT 31.730 0.300 32.070 0.985 ;
        RECT 34.025 0.300 34.255 1.050 ;
        RECT 0.000 -0.300 34.720 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 2.760 1.595 3.390 ;
        RECT 3.505 2.760 3.735 3.390 ;
        RECT 5.745 2.760 5.975 3.390 ;
        RECT 7.985 2.820 8.215 3.390 ;
        RECT 10.325 2.820 10.555 3.390 ;
        RECT 7.985 2.760 10.555 2.820 ;
        RECT 1.365 2.530 10.555 2.760 ;
        RECT 10.325 1.995 10.555 2.530 ;
        RECT 10.325 1.765 21.280 1.995 ;
        RECT 23.860 1.765 32.660 1.995 ;
        RECT 10.325 1.505 10.555 1.765 ;
        RECT 1.365 1.270 10.555 1.505 ;
        RECT 1.365 0.685 1.595 1.270 ;
        RECT 3.605 0.685 3.835 1.270 ;
        RECT 5.845 0.685 6.075 1.270 ;
        RECT 8.085 0.685 8.315 1.270 ;
        RECT 10.325 0.685 10.555 1.270 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__clkbuf_20
MACRO gf180mcu_fd_sc_mcu7t5v0__clkinv_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkinv_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.898000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 0.970 1.030 2.950 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.748000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.260 0.600 1.595 3.370 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 2.240 4.220 ;
        RECT 0.245 2.480 0.475 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 2.670 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.040 ;
        RECT 0.000 -0.300 2.240 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__clkinv_1
MACRO gf180mcu_fd_sc_mcu7t5v0__clkinv_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkinv_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.796000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 2.120 1.035 2.875 ;
        RECT 0.705 1.735 1.970 2.120 ;
        RECT 0.705 1.190 1.035 1.735 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.006000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 2.735 1.495 3.380 ;
        RECT 1.265 2.360 2.710 2.735 ;
        RECT 2.330 1.505 2.710 2.360 ;
        RECT 1.365 1.270 2.710 1.505 ;
        RECT 1.365 0.680 1.595 1.270 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 3.360 4.220 ;
        RECT 0.245 2.530 0.475 3.620 ;
        RECT 2.330 2.965 2.670 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 3.790 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 3.790 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.040 ;
        RECT 2.485 0.300 2.715 1.040 ;
        RECT 0.000 -0.300 3.360 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__clkinv_2
MACRO gf180mcu_fd_sc_mcu7t5v0__clkinv_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkinv_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.694000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 1.740 2.855 2.120 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.754000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 2.735 1.495 3.380 ;
        RECT 3.450 2.735 3.835 3.380 ;
        RECT 1.265 2.360 3.835 2.735 ;
        RECT 3.460 1.505 3.835 2.360 ;
        RECT 1.365 1.270 3.835 1.505 ;
        RECT 1.365 0.700 1.595 1.270 ;
        RECT 3.450 0.650 3.835 1.270 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 4.480 4.220 ;
        RECT 0.245 2.550 0.475 3.620 ;
        RECT 2.330 2.965 2.670 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 4.910 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.040 ;
        RECT 2.485 0.300 2.715 1.040 ;
        RECT 0.000 -0.300 4.480 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__clkinv_3
MACRO gf180mcu_fd_sc_mcu7t5v0__clkinv_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkinv_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.592000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 1.765 2.710 2.150 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.256000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 2.705 1.595 3.270 ;
        RECT 3.450 2.705 3.835 3.270 ;
        RECT 1.365 2.385 3.835 2.705 ;
        RECT 3.450 1.535 3.835 2.385 ;
        RECT 1.365 1.215 3.835 1.535 ;
        RECT 1.365 0.700 1.595 1.215 ;
        RECT 3.450 0.700 3.835 1.215 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.600 4.220 ;
        RECT 0.245 2.590 0.475 3.620 ;
        RECT 2.430 2.965 2.770 3.620 ;
        RECT 4.725 2.590 4.955 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 6.030 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.040 ;
        RECT 2.430 0.300 2.770 0.985 ;
        RECT 4.725 0.300 4.955 1.040 ;
        RECT 0.000 -0.300 5.600 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__clkinv_4
MACRO gf180mcu_fd_sc_mcu7t5v0__clkinv_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkinv_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 7.184000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 1.765 3.790 2.150 ;
        RECT 5.330 1.765 8.960 2.150 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.024000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 2.730 1.495 3.380 ;
        RECT 3.505 2.730 3.735 3.380 ;
        RECT 1.265 2.725 3.735 2.730 ;
        RECT 5.745 2.725 5.975 3.380 ;
        RECT 7.985 2.725 8.215 3.380 ;
        RECT 1.265 2.410 8.215 2.725 ;
        RECT 4.570 1.535 4.950 2.410 ;
        RECT 1.365 1.215 8.315 1.535 ;
        RECT 1.365 0.700 1.595 1.215 ;
        RECT 3.605 0.700 3.835 1.215 ;
        RECT 5.845 0.700 6.075 1.215 ;
        RECT 8.085 0.700 8.315 1.215 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 10.080 4.220 ;
        RECT 0.245 2.550 0.475 3.620 ;
        RECT 2.330 2.965 2.670 3.620 ;
        RECT 4.570 2.965 4.910 3.620 ;
        RECT 6.810 2.965 7.150 3.620 ;
        RECT 9.105 2.550 9.335 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 10.510 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.040 ;
        RECT 2.430 0.300 2.770 0.985 ;
        RECT 4.670 0.300 5.010 0.985 ;
        RECT 6.910 0.300 7.250 0.985 ;
        RECT 9.205 0.300 9.435 1.040 ;
        RECT 0.000 -0.300 10.080 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__clkinv_8
MACRO gf180mcu_fd_sc_mcu7t5v0__clkinv_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkinv_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 10.776000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.620 1.765 5.820 2.150 ;
        RECT 7.990 1.765 13.540 2.150 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.036000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 3.050 1.495 3.380 ;
        RECT 3.505 3.050 3.735 3.380 ;
        RECT 5.690 3.050 6.070 3.380 ;
        RECT 1.265 3.045 6.070 3.050 ;
        RECT 7.985 3.045 8.215 3.380 ;
        RECT 10.225 3.045 10.455 3.380 ;
        RECT 12.465 3.045 12.695 3.380 ;
        RECT 1.265 2.570 12.695 3.045 ;
        RECT 6.550 1.535 7.450 2.570 ;
        RECT 1.365 1.100 12.795 1.535 ;
        RECT 1.365 0.585 1.595 1.100 ;
        RECT 3.605 0.585 3.835 1.100 ;
        RECT 5.845 0.585 6.075 1.100 ;
        RECT 8.085 0.585 8.315 1.100 ;
        RECT 10.325 0.585 10.555 1.100 ;
        RECT 12.565 0.585 12.795 1.100 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 14.560 4.220 ;
        RECT 0.245 2.570 0.475 3.620 ;
        RECT 2.330 3.280 2.670 3.620 ;
        RECT 4.570 3.280 4.910 3.620 ;
        RECT 6.810 3.280 7.150 3.620 ;
        RECT 9.050 3.280 9.390 3.620 ;
        RECT 11.290 3.280 11.630 3.620 ;
        RECT 13.585 2.570 13.815 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 14.990 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 0.925 ;
        RECT 2.430 0.300 2.770 0.870 ;
        RECT 4.670 0.300 5.010 0.870 ;
        RECT 6.910 0.300 7.250 0.870 ;
        RECT 9.150 0.300 9.490 0.870 ;
        RECT 11.390 0.300 11.730 0.870 ;
        RECT 13.685 0.300 13.915 0.925 ;
        RECT 0.000 -0.300 14.560 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__clkinv_12
MACRO gf180mcu_fd_sc_mcu7t5v0__clkinv_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkinv_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.040 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 14.368000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.640 1.760 8.130 2.150 ;
        RECT 10.280 1.765 17.670 2.150 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 8.047999 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 3.055 1.495 3.380 ;
        RECT 3.505 3.055 3.735 3.380 ;
        RECT 5.745 3.055 5.975 3.380 ;
        RECT 7.930 3.055 8.310 3.380 ;
        RECT 10.225 3.055 10.455 3.380 ;
        RECT 12.465 3.055 12.695 3.380 ;
        RECT 14.705 3.055 14.935 3.380 ;
        RECT 16.945 3.055 17.175 3.380 ;
        RECT 1.265 2.475 17.175 3.055 ;
        RECT 8.790 1.455 9.690 2.475 ;
        RECT 1.310 0.875 17.330 1.455 ;
        RECT 1.310 0.530 1.650 0.875 ;
        RECT 3.550 0.530 3.890 0.875 ;
        RECT 5.790 0.530 6.130 0.875 ;
        RECT 8.030 0.530 8.370 0.875 ;
        RECT 10.270 0.530 10.610 0.875 ;
        RECT 12.510 0.530 12.850 0.875 ;
        RECT 14.750 0.530 15.090 0.875 ;
        RECT 16.990 0.530 17.330 0.875 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 19.040 4.220 ;
        RECT 0.245 2.570 0.475 3.620 ;
        RECT 2.330 3.285 2.670 3.620 ;
        RECT 4.570 3.285 4.910 3.620 ;
        RECT 6.810 3.285 7.150 3.620 ;
        RECT 9.050 3.285 9.390 3.620 ;
        RECT 11.290 3.285 11.630 3.620 ;
        RECT 13.530 3.285 13.870 3.620 ;
        RECT 15.770 3.285 16.110 3.620 ;
        RECT 18.065 2.530 18.295 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 19.470 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 19.470 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 0.700 ;
        RECT 2.430 0.300 2.770 0.645 ;
        RECT 4.670 0.300 5.010 0.645 ;
        RECT 6.910 0.300 7.250 0.645 ;
        RECT 9.150 0.300 9.490 0.645 ;
        RECT 11.390 0.300 11.730 0.645 ;
        RECT 13.630 0.300 13.970 0.645 ;
        RECT 15.870 0.300 16.210 0.645 ;
        RECT 18.165 0.300 18.395 0.700 ;
        RECT 0.000 -0.300 19.040 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__clkinv_16
MACRO gf180mcu_fd_sc_mcu7t5v0__clkinv_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkinv_20 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.520 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 17.959999 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 1.740 9.900 2.120 ;
        RECT 12.520 1.740 22.400 2.120 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 10.059999 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.055 1.595 3.380 ;
        RECT 3.505 3.055 3.735 3.380 ;
        RECT 5.745 3.055 5.975 3.380 ;
        RECT 7.985 3.055 8.215 3.380 ;
        RECT 10.170 3.055 10.550 3.380 ;
        RECT 12.465 3.055 12.695 3.380 ;
        RECT 14.705 3.055 14.935 3.380 ;
        RECT 16.945 3.055 17.175 3.380 ;
        RECT 19.185 3.055 19.415 3.380 ;
        RECT 21.425 3.055 21.655 3.380 ;
        RECT 1.365 2.350 21.655 3.055 ;
        RECT 11.030 1.505 11.930 2.350 ;
        RECT 1.310 0.875 21.810 1.505 ;
        RECT 1.310 0.535 1.650 0.875 ;
        RECT 3.550 0.535 3.890 0.875 ;
        RECT 5.790 0.535 6.130 0.875 ;
        RECT 8.030 0.535 8.370 0.875 ;
        RECT 10.270 0.535 10.610 0.875 ;
        RECT 12.510 0.535 12.850 0.875 ;
        RECT 14.750 0.535 15.090 0.875 ;
        RECT 16.990 0.535 17.330 0.875 ;
        RECT 19.230 0.535 19.570 0.875 ;
        RECT 21.470 0.535 21.810 0.875 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 23.520 4.220 ;
        RECT 0.245 2.530 0.475 3.620 ;
        RECT 2.330 3.285 2.670 3.620 ;
        RECT 4.570 3.285 4.910 3.620 ;
        RECT 6.810 3.285 7.150 3.620 ;
        RECT 9.050 3.285 9.390 3.620 ;
        RECT 11.290 3.285 11.630 3.620 ;
        RECT 13.530 3.285 13.870 3.620 ;
        RECT 15.770 3.285 16.110 3.620 ;
        RECT 18.010 3.285 18.350 3.620 ;
        RECT 20.250 3.285 20.590 3.620 ;
        RECT 22.545 2.530 22.775 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 23.950 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 23.950 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 0.700 ;
        RECT 2.430 0.300 2.770 0.645 ;
        RECT 4.670 0.300 5.010 0.645 ;
        RECT 6.910 0.300 7.250 0.645 ;
        RECT 9.150 0.300 9.490 0.645 ;
        RECT 11.390 0.300 11.730 0.645 ;
        RECT 13.630 0.300 13.970 0.645 ;
        RECT 15.870 0.300 16.210 0.645 ;
        RECT 18.110 0.300 18.450 0.645 ;
        RECT 20.350 0.300 20.690 0.645 ;
        RECT 22.590 0.300 22.930 0.645 ;
        RECT 0.000 -0.300 23.520 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__clkinv_20
MACRO gf180mcu_fd_sc_mcu7t5v0__dffnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.800 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.463500 ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 1.770 4.390 2.150 ;
    END
  END D
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.711500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.280 1.770 1.590 2.130 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.858000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.770 0.810 16.350 2.985 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 16.800 4.220 ;
        RECT 1.440 2.930 1.780 3.620 ;
        RECT 3.180 3.005 3.520 3.620 ;
        RECT 7.705 2.700 8.045 3.620 ;
        RECT 12.850 3.280 13.190 3.620 ;
        RECT 14.845 2.755 15.185 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 17.230 4.350 ;
        RECT -0.430 1.760 7.265 1.885 ;
        RECT 14.620 1.760 17.230 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 7.265 1.760 14.620 1.885 ;
        RECT -0.430 -0.430 17.230 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.440 0.300 1.780 0.915 ;
        RECT 3.280 0.300 3.620 1.075 ;
        RECT 7.700 0.300 8.040 0.810 ;
        RECT 12.720 0.300 13.060 0.950 ;
        RECT 15.000 0.300 15.230 0.690 ;
        RECT 0.000 -0.300 16.800 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.475 2.590 0.705 3.225 ;
        RECT 2.515 2.710 2.845 3.225 ;
        RECT 3.830 3.160 6.355 3.390 ;
        RECT 3.830 2.710 4.060 3.160 ;
        RECT 13.430 3.100 14.615 3.330 ;
        RECT 13.430 3.050 13.660 3.100 ;
        RECT 0.475 2.360 2.165 2.590 ;
        RECT 1.935 1.375 2.165 2.360 ;
        RECT 0.375 1.145 2.165 1.375 ;
        RECT 2.515 2.480 4.060 2.710 ;
        RECT 4.420 2.645 5.290 2.875 ;
        RECT 0.375 0.735 0.605 1.145 ;
        RECT 2.515 0.735 2.845 2.480 ;
        RECT 5.055 1.075 5.290 2.645 ;
        RECT 4.400 0.845 5.290 1.075 ;
        RECT 5.575 2.050 5.915 2.795 ;
        RECT 9.040 2.390 9.380 2.930 ;
        RECT 7.095 2.050 9.380 2.390 ;
        RECT 5.575 1.820 6.780 2.050 ;
        RECT 5.575 0.790 5.805 1.820 ;
        RECT 6.550 1.730 6.780 1.820 ;
        RECT 6.090 1.270 6.320 1.590 ;
        RECT 6.550 1.500 8.700 1.730 ;
        RECT 6.090 1.040 8.560 1.270 ;
        RECT 8.330 0.760 8.560 1.040 ;
        RECT 9.040 0.990 9.380 2.050 ;
        RECT 10.160 2.585 10.500 2.930 ;
        RECT 11.790 2.815 13.660 3.050 ;
        RECT 10.160 2.355 13.630 2.585 ;
        RECT 10.160 0.990 10.500 2.355 ;
        RECT 13.290 2.105 13.630 2.355 ;
        RECT 11.195 0.760 11.425 2.095 ;
        RECT 13.925 1.885 14.155 2.850 ;
        RECT 14.385 2.345 14.615 3.100 ;
        RECT 14.385 2.115 15.460 2.345 ;
        RECT 13.925 1.875 15.000 1.885 ;
        RECT 12.175 1.640 15.000 1.875 ;
        RECT 13.900 1.500 15.000 1.640 ;
        RECT 11.655 1.180 13.520 1.410 ;
        RECT 11.655 0.890 11.885 1.180 ;
        RECT 8.330 0.530 11.425 0.760 ;
        RECT 13.290 0.760 13.520 1.180 ;
        RECT 13.900 0.990 14.240 1.500 ;
        RECT 15.230 1.150 15.460 2.115 ;
        RECT 14.540 0.920 15.460 1.150 ;
        RECT 14.540 0.760 14.770 0.920 ;
        RECT 13.290 0.530 14.770 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnq_1
MACRO gf180mcu_fd_sc_mcu7t5v0__dffnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.480 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.463500 ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 1.770 4.390 2.150 ;
    END
  END D
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.711500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.280 1.770 1.590 2.130 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.401600 ;
    PORT
      LAYER Metal1 ;
        RECT 15.965 2.150 16.315 2.930 ;
        RECT 15.965 1.770 17.270 2.150 ;
        RECT 16.285 0.990 16.625 1.770 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 18.480 4.220 ;
        RECT 1.440 2.930 1.780 3.620 ;
        RECT 3.180 3.005 3.520 3.620 ;
        RECT 7.705 2.700 8.045 3.620 ;
        RECT 12.850 3.280 13.190 3.620 ;
        RECT 14.845 2.815 15.185 3.620 ;
        RECT 17.040 2.760 17.270 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 18.910 4.350 ;
        RECT -0.430 1.760 7.265 1.885 ;
        RECT 17.275 1.760 18.910 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 7.265 1.760 17.275 1.885 ;
        RECT -0.430 -0.430 18.910 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.440 0.300 1.780 0.915 ;
        RECT 3.280 0.300 3.620 1.075 ;
        RECT 7.700 0.300 8.040 0.810 ;
        RECT 12.850 0.300 13.190 0.635 ;
        RECT 15.000 0.300 15.230 0.690 ;
        RECT 17.625 0.300 17.965 0.635 ;
        RECT 0.000 -0.300 18.480 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.475 2.590 0.705 3.225 ;
        RECT 2.515 2.710 2.845 3.225 ;
        RECT 3.830 3.160 6.355 3.390 ;
        RECT 3.830 2.710 4.060 3.160 ;
        RECT 13.430 3.100 14.615 3.330 ;
        RECT 13.430 3.050 13.660 3.100 ;
        RECT 0.475 2.360 2.165 2.590 ;
        RECT 1.935 1.375 2.165 2.360 ;
        RECT 0.375 1.145 2.165 1.375 ;
        RECT 2.515 2.480 4.060 2.710 ;
        RECT 4.420 2.645 5.290 2.875 ;
        RECT 0.375 0.735 0.605 1.145 ;
        RECT 2.515 0.735 2.845 2.480 ;
        RECT 5.055 1.075 5.290 2.645 ;
        RECT 4.400 0.845 5.290 1.075 ;
        RECT 5.575 2.050 5.915 2.795 ;
        RECT 9.040 2.390 9.380 2.930 ;
        RECT 7.095 2.050 9.380 2.390 ;
        RECT 5.575 1.820 6.780 2.050 ;
        RECT 5.575 0.790 5.805 1.820 ;
        RECT 6.550 1.730 6.780 1.820 ;
        RECT 6.090 1.270 6.320 1.590 ;
        RECT 6.550 1.500 8.700 1.730 ;
        RECT 6.090 1.040 8.560 1.270 ;
        RECT 8.330 0.760 8.560 1.040 ;
        RECT 9.040 0.990 9.380 2.050 ;
        RECT 10.160 2.585 10.500 2.930 ;
        RECT 11.790 2.815 13.660 3.050 ;
        RECT 10.160 2.355 13.575 2.585 ;
        RECT 10.160 0.990 10.500 2.355 ;
        RECT 13.345 2.050 13.575 2.355 ;
        RECT 13.925 2.055 14.155 2.850 ;
        RECT 14.385 2.515 14.615 3.100 ;
        RECT 14.385 2.285 15.645 2.515 ;
        RECT 11.170 0.760 11.510 2.040 ;
        RECT 13.925 1.730 15.075 2.055 ;
        RECT 12.410 1.715 15.075 1.730 ;
        RECT 12.410 1.495 14.310 1.715 ;
        RECT 8.330 0.530 11.510 0.760 ;
        RECT 11.745 0.865 13.650 1.095 ;
        RECT 13.970 0.990 14.310 1.495 ;
        RECT 15.415 1.150 15.645 2.285 ;
        RECT 11.745 0.675 11.975 0.865 ;
        RECT 13.420 0.760 13.650 0.865 ;
        RECT 14.540 0.920 15.645 1.150 ;
        RECT 14.540 0.760 14.770 0.920 ;
        RECT 13.420 0.530 14.770 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnq_2
MACRO gf180mcu_fd_sc_mcu7t5v0__dffnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.463500 ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 1.770 4.390 2.150 ;
    END
  END D
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.711500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.280 1.770 1.590 2.130 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.525900 ;
    PORT
      LAYER Metal1 ;
        RECT 16.490 2.595 16.840 2.930 ;
        RECT 18.870 2.595 19.510 2.930 ;
        RECT 16.490 2.245 19.510 2.595 ;
        RECT 18.570 1.555 19.510 2.245 ;
        RECT 16.490 1.325 19.510 1.555 ;
        RECT 16.490 0.990 16.830 1.325 ;
        RECT 19.170 0.990 19.510 1.325 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 21.280 4.220 ;
        RECT 1.440 2.930 1.780 3.620 ;
        RECT 3.180 3.005 3.520 3.620 ;
        RECT 7.705 2.700 8.045 3.620 ;
        RECT 12.850 3.280 13.190 3.620 ;
        RECT 15.250 2.815 15.590 3.620 ;
        RECT 17.730 3.285 18.070 3.620 ;
        RECT 20.510 2.815 20.850 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 21.710 4.350 ;
        RECT -0.430 1.760 7.265 1.885 ;
        RECT 20.350 1.760 21.710 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 7.265 1.760 20.350 1.885 ;
        RECT -0.430 -0.430 21.710 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.440 0.300 1.780 0.915 ;
        RECT 3.280 0.300 3.620 1.075 ;
        RECT 7.700 0.300 8.040 0.810 ;
        RECT 12.850 0.300 13.190 0.635 ;
        RECT 15.205 0.300 15.435 0.690 ;
        RECT 17.830 0.300 18.170 0.635 ;
        RECT 20.565 0.300 20.795 0.765 ;
        RECT 0.000 -0.300 21.280 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.475 2.590 0.705 3.225 ;
        RECT 2.515 2.710 2.845 3.225 ;
        RECT 3.830 3.160 6.355 3.390 ;
        RECT 3.830 2.710 4.060 3.160 ;
        RECT 13.500 3.050 15.020 3.255 ;
        RECT 11.790 3.025 15.020 3.050 ;
        RECT 0.475 2.360 2.165 2.590 ;
        RECT 1.935 1.375 2.165 2.360 ;
        RECT 0.375 1.145 2.165 1.375 ;
        RECT 2.515 2.480 4.060 2.710 ;
        RECT 4.420 2.645 5.290 2.875 ;
        RECT 0.375 0.735 0.605 1.145 ;
        RECT 2.515 0.735 2.845 2.480 ;
        RECT 5.055 1.075 5.290 2.645 ;
        RECT 4.400 0.845 5.290 1.075 ;
        RECT 5.575 2.050 5.915 2.795 ;
        RECT 9.040 2.390 9.380 2.930 ;
        RECT 7.095 2.050 9.380 2.390 ;
        RECT 5.575 1.820 6.780 2.050 ;
        RECT 5.575 0.790 5.805 1.820 ;
        RECT 6.550 1.730 6.780 1.820 ;
        RECT 6.090 1.270 6.320 1.590 ;
        RECT 6.550 1.500 8.700 1.730 ;
        RECT 6.090 1.040 8.560 1.270 ;
        RECT 8.330 0.760 8.560 1.040 ;
        RECT 9.040 0.990 9.380 2.050 ;
        RECT 10.160 2.585 10.500 2.930 ;
        RECT 11.790 2.815 13.730 3.025 ;
        RECT 10.160 2.355 13.770 2.585 ;
        RECT 10.160 0.990 10.500 2.355 ;
        RECT 13.430 2.105 13.770 2.355 ;
        RECT 11.170 0.760 11.510 2.040 ;
        RECT 14.090 2.015 14.430 2.795 ;
        RECT 14.790 2.525 15.020 3.025 ;
        RECT 15.825 3.160 17.500 3.390 ;
        RECT 15.825 2.525 16.055 3.160 ;
        RECT 17.270 3.055 17.500 3.160 ;
        RECT 18.300 3.160 20.130 3.390 ;
        RECT 18.300 3.055 18.530 3.160 ;
        RECT 17.270 2.825 18.530 3.055 ;
        RECT 14.790 2.295 16.055 2.525 ;
        RECT 14.090 1.785 17.910 2.015 ;
        RECT 14.090 1.730 14.490 1.785 ;
        RECT 12.410 1.495 14.490 1.730 ;
        RECT 8.330 0.530 11.510 0.760 ;
        RECT 11.745 0.865 13.650 1.095 ;
        RECT 14.150 0.990 14.490 1.495 ;
        RECT 11.745 0.675 11.975 0.865 ;
        RECT 13.420 0.760 13.650 0.865 ;
        RECT 14.745 0.920 15.895 1.150 ;
        RECT 14.745 0.760 14.975 0.920 ;
        RECT 13.420 0.530 14.975 0.760 ;
        RECT 15.665 0.760 15.895 0.920 ;
        RECT 17.370 0.865 18.630 1.095 ;
        RECT 17.370 0.760 17.600 0.865 ;
        RECT 15.665 0.530 17.600 0.760 ;
        RECT 18.400 0.760 18.630 0.865 ;
        RECT 19.900 0.760 20.130 3.160 ;
        RECT 18.400 0.530 20.130 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnq_4
MACRO gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.040 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.614000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.890 1.770 3.895 2.150 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.318000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.650 1.020 15.140 1.830 ;
        RECT 14.650 0.600 16.300 1.020 ;
    END
  END RN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.675500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.290 1.770 1.575 2.150 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.866800 ;
    PORT
      LAYER Metal1 ;
        RECT 18.365 2.765 18.920 3.320 ;
        RECT 17.450 2.330 18.920 2.765 ;
        RECT 18.570 0.830 18.920 2.330 ;
        RECT 18.380 0.600 18.920 0.830 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 19.040 4.220 ;
        RECT 1.310 2.930 1.650 3.620 ;
        RECT 3.170 2.845 3.510 3.620 ;
        RECT 7.590 3.005 7.930 3.620 ;
        RECT 9.605 2.790 9.835 3.620 ;
        RECT 14.220 3.280 14.560 3.620 ;
        RECT 16.595 2.690 16.825 3.620 ;
        RECT 17.415 3.160 17.645 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 19.470 4.350 ;
        RECT -0.430 1.770 9.525 1.885 ;
        RECT -0.430 1.760 2.960 1.770 ;
        RECT 17.040 1.760 19.470 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 9.525 1.770 17.040 1.885 ;
        RECT 2.960 1.760 17.040 1.770 ;
        RECT -0.430 -0.430 19.470 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.915 ;
        RECT 3.150 0.300 3.490 1.075 ;
        RECT 8.530 0.300 8.870 0.915 ;
        RECT 14.175 0.300 14.405 1.130 ;
        RECT 17.315 0.300 17.545 0.930 ;
        RECT 0.000 -0.300 19.040 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.785 3.160 5.015 3.390 ;
        RECT 0.345 2.700 0.575 2.805 ;
        RECT 0.345 2.465 2.035 2.700 ;
        RECT 1.805 1.375 2.035 2.465 ;
        RECT 0.245 1.145 2.035 1.375 ;
        RECT 2.385 2.610 2.615 2.805 ;
        RECT 3.785 2.610 4.015 3.160 ;
        RECT 2.385 2.380 4.015 2.610 ;
        RECT 0.245 0.630 0.475 1.145 ;
        RECT 2.385 0.970 2.615 2.380 ;
        RECT 2.385 0.630 2.715 0.970 ;
        RECT 4.245 0.790 4.555 2.800 ;
        RECT 4.785 1.555 5.015 3.160 ;
        RECT 11.875 3.160 13.900 3.390 ;
        RECT 5.265 2.315 5.495 2.800 ;
        RECT 6.285 2.775 6.515 3.115 ;
        RECT 8.160 2.830 9.170 3.060 ;
        RECT 8.160 2.775 8.390 2.830 ;
        RECT 6.285 2.545 8.390 2.775 ;
        RECT 8.620 2.315 10.330 2.470 ;
        RECT 5.265 2.240 10.330 2.315 ;
        RECT 5.265 2.085 8.850 2.240 ;
        RECT 5.265 0.790 5.675 2.085 ;
        RECT 10.625 2.010 10.855 3.130 ;
        RECT 11.875 2.405 12.105 3.160 ;
        RECT 13.670 3.050 13.900 3.160 ;
        RECT 14.790 3.160 16.365 3.390 ;
        RECT 14.790 3.050 15.020 3.160 ;
        RECT 10.060 1.855 10.855 2.010 ;
        RECT 6.930 1.780 10.855 1.855 ;
        RECT 11.645 2.065 12.105 2.405 ;
        RECT 6.930 1.625 10.430 1.780 ;
        RECT 6.170 1.395 6.515 1.565 ;
        RECT 6.170 1.165 9.330 1.395 ;
        RECT 9.100 0.760 9.330 1.165 ;
        RECT 10.090 0.990 10.430 1.625 ;
        RECT 11.025 0.760 11.255 1.620 ;
        RECT 11.645 0.990 11.995 2.065 ;
        RECT 12.395 0.760 12.625 2.525 ;
        RECT 12.980 0.820 13.320 2.930 ;
        RECT 13.670 2.815 15.020 3.050 ;
        RECT 15.450 2.470 15.790 2.930 ;
        RECT 13.560 2.235 15.790 2.470 ;
        RECT 15.560 1.735 15.790 2.235 ;
        RECT 16.135 2.375 16.365 3.160 ;
        RECT 16.135 2.035 16.385 2.375 ;
        RECT 15.560 1.505 18.040 1.735 ;
        RECT 16.595 0.790 16.825 1.505 ;
        RECT 9.100 0.530 12.625 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
MACRO gf180mcu_fd_sc_mcu7t5v0__dffnrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnrnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.160 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.614000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.890 1.770 3.895 2.150 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.393000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.650 0.650 15.140 1.590 ;
    END
  END RN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.675500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 1.575 2.150 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.029600 ;
    PORT
      LAYER Metal1 ;
        RECT 18.380 2.765 18.720 3.235 ;
        RECT 18.380 2.330 19.510 2.765 ;
        RECT 19.130 1.175 19.510 2.330 ;
        RECT 18.435 0.945 19.510 1.175 ;
        RECT 18.435 0.790 18.665 0.945 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 20.160 4.220 ;
        RECT 1.310 2.930 1.650 3.620 ;
        RECT 3.170 2.845 3.510 3.620 ;
        RECT 7.590 3.005 7.930 3.620 ;
        RECT 9.605 2.790 9.835 3.620 ;
        RECT 14.220 3.280 14.560 3.620 ;
        RECT 16.595 2.690 16.825 3.620 ;
        RECT 17.415 2.690 17.645 3.620 ;
        RECT 19.455 3.160 19.685 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 20.590 4.350 ;
        RECT -0.430 1.770 9.525 1.885 ;
        RECT -0.430 1.760 2.960 1.770 ;
        RECT 17.020 1.760 20.590 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 9.525 1.770 17.020 1.885 ;
        RECT 2.960 1.760 17.020 1.770 ;
        RECT -0.430 -0.430 20.590 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.915 ;
        RECT 3.150 0.300 3.490 1.075 ;
        RECT 8.530 0.300 8.870 0.915 ;
        RECT 14.175 0.300 14.405 1.130 ;
        RECT 17.315 0.300 17.545 0.765 ;
        RECT 19.500 0.300 19.840 0.715 ;
        RECT 0.000 -0.300 20.160 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.785 3.160 5.015 3.390 ;
        RECT 0.345 2.700 0.575 2.805 ;
        RECT 0.345 2.465 2.035 2.700 ;
        RECT 1.805 1.375 2.035 2.465 ;
        RECT 0.245 1.145 2.035 1.375 ;
        RECT 2.385 2.610 2.615 2.805 ;
        RECT 3.785 2.610 4.015 3.160 ;
        RECT 2.385 2.380 4.015 2.610 ;
        RECT 0.245 0.630 0.475 1.145 ;
        RECT 2.385 0.970 2.615 2.380 ;
        RECT 2.385 0.630 2.715 0.970 ;
        RECT 4.245 0.790 4.555 2.800 ;
        RECT 4.785 1.555 5.015 3.160 ;
        RECT 11.875 3.160 13.900 3.390 ;
        RECT 5.265 2.315 5.495 2.800 ;
        RECT 6.285 2.775 6.515 3.115 ;
        RECT 8.160 2.830 9.170 3.060 ;
        RECT 8.160 2.775 8.390 2.830 ;
        RECT 6.285 2.545 8.390 2.775 ;
        RECT 8.620 2.315 10.330 2.470 ;
        RECT 5.265 2.240 10.330 2.315 ;
        RECT 5.265 2.085 8.850 2.240 ;
        RECT 5.265 0.790 5.675 2.085 ;
        RECT 10.625 2.010 10.855 3.130 ;
        RECT 11.875 2.405 12.105 3.160 ;
        RECT 13.670 3.050 13.900 3.160 ;
        RECT 14.790 3.155 16.365 3.390 ;
        RECT 14.790 3.050 15.020 3.155 ;
        RECT 10.060 1.855 10.855 2.010 ;
        RECT 6.930 1.780 10.855 1.855 ;
        RECT 11.645 2.065 12.105 2.405 ;
        RECT 6.930 1.625 10.430 1.780 ;
        RECT 6.170 1.395 6.515 1.565 ;
        RECT 6.170 1.165 9.330 1.395 ;
        RECT 9.100 0.760 9.330 1.165 ;
        RECT 10.090 0.990 10.430 1.625 ;
        RECT 11.025 0.760 11.255 1.620 ;
        RECT 11.645 0.990 11.995 2.065 ;
        RECT 12.395 0.760 12.625 2.525 ;
        RECT 12.980 0.820 13.320 2.930 ;
        RECT 13.670 2.815 15.020 3.050 ;
        RECT 15.450 2.470 15.790 2.870 ;
        RECT 13.560 2.235 15.790 2.470 ;
        RECT 13.560 1.770 13.900 2.235 ;
        RECT 15.560 1.735 15.790 2.235 ;
        RECT 16.135 2.375 16.365 3.155 ;
        RECT 16.135 2.035 16.385 2.375 ;
        RECT 15.560 1.505 18.610 1.735 ;
        RECT 9.100 0.530 12.625 0.760 ;
        RECT 16.595 0.740 16.825 1.505 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnrnq_2
MACRO gf180mcu_fd_sc_mcu7t5v0__dffnrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnrnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.400 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.614000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.890 1.770 3.895 2.150 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.395500 ;
    PORT
      LAYER Metal1 ;
        RECT 14.650 0.650 15.140 1.590 ;
    END
  END RN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.675500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.770 1.575 2.150 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.080000 ;
    PORT
      LAYER Metal1 ;
        RECT 18.380 2.765 18.720 3.235 ;
        RECT 20.420 2.765 20.760 3.235 ;
        RECT 18.380 2.330 21.190 2.765 ;
        RECT 20.810 1.175 21.190 2.330 ;
        RECT 18.435 0.945 21.190 1.175 ;
        RECT 18.435 0.790 18.665 0.945 ;
        RECT 20.635 0.790 21.190 0.945 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 22.400 4.220 ;
        RECT 1.310 2.930 1.650 3.620 ;
        RECT 3.170 2.845 3.510 3.620 ;
        RECT 7.590 3.005 7.930 3.620 ;
        RECT 9.605 2.790 9.835 3.620 ;
        RECT 14.220 3.280 14.560 3.620 ;
        RECT 16.595 2.690 16.825 3.620 ;
        RECT 17.415 2.690 17.645 3.620 ;
        RECT 19.455 3.160 19.685 3.620 ;
        RECT 21.495 2.690 21.725 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 22.830 4.350 ;
        RECT -0.430 1.770 9.525 1.885 ;
        RECT -0.430 1.760 2.960 1.770 ;
        RECT 17.000 1.760 22.830 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 9.525 1.770 17.000 1.885 ;
        RECT 2.960 1.760 17.000 1.770 ;
        RECT -0.430 -0.430 22.830 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.915 ;
        RECT 3.150 0.300 3.490 1.075 ;
        RECT 8.530 0.300 8.870 0.915 ;
        RECT 14.175 0.300 14.405 1.130 ;
        RECT 17.315 0.300 17.545 0.765 ;
        RECT 19.500 0.300 19.840 0.715 ;
        RECT 21.795 0.300 22.025 0.765 ;
        RECT 0.000 -0.300 22.400 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.785 3.160 5.015 3.390 ;
        RECT 0.345 2.700 0.575 2.805 ;
        RECT 0.345 2.465 2.035 2.700 ;
        RECT 1.805 1.375 2.035 2.465 ;
        RECT 0.245 1.145 2.035 1.375 ;
        RECT 2.385 2.610 2.615 2.805 ;
        RECT 3.785 2.610 4.015 3.160 ;
        RECT 2.385 2.380 4.015 2.610 ;
        RECT 0.245 0.630 0.475 1.145 ;
        RECT 2.385 0.970 2.615 2.380 ;
        RECT 2.385 0.630 2.715 0.970 ;
        RECT 4.245 0.790 4.555 2.800 ;
        RECT 4.785 1.555 5.015 3.160 ;
        RECT 11.875 3.160 13.900 3.390 ;
        RECT 5.265 2.315 5.495 2.800 ;
        RECT 6.285 2.775 6.515 3.115 ;
        RECT 8.160 2.830 9.170 3.060 ;
        RECT 8.160 2.775 8.390 2.830 ;
        RECT 6.285 2.545 8.390 2.775 ;
        RECT 8.620 2.315 10.330 2.470 ;
        RECT 5.265 2.240 10.330 2.315 ;
        RECT 5.265 2.085 8.850 2.240 ;
        RECT 5.265 0.790 5.675 2.085 ;
        RECT 10.625 2.010 10.855 3.130 ;
        RECT 11.875 2.405 12.105 3.160 ;
        RECT 13.670 3.050 13.900 3.160 ;
        RECT 14.790 3.155 16.365 3.390 ;
        RECT 14.790 3.050 15.020 3.155 ;
        RECT 10.060 1.855 10.855 2.010 ;
        RECT 6.930 1.780 10.855 1.855 ;
        RECT 11.645 2.065 12.105 2.405 ;
        RECT 6.930 1.625 10.430 1.780 ;
        RECT 6.170 1.395 6.515 1.565 ;
        RECT 6.170 1.165 9.330 1.395 ;
        RECT 9.100 0.760 9.330 1.165 ;
        RECT 10.090 0.990 10.430 1.625 ;
        RECT 11.025 0.760 11.255 1.620 ;
        RECT 11.645 0.990 11.995 2.065 ;
        RECT 12.395 0.760 12.625 2.525 ;
        RECT 12.980 0.820 13.320 2.930 ;
        RECT 13.670 2.815 15.020 3.050 ;
        RECT 15.450 2.470 15.790 2.870 ;
        RECT 13.560 2.235 15.790 2.470 ;
        RECT 13.560 1.770 13.900 2.235 ;
        RECT 15.560 1.665 15.790 2.235 ;
        RECT 16.135 2.375 16.365 3.155 ;
        RECT 16.135 2.035 16.385 2.375 ;
        RECT 15.560 1.435 20.280 1.665 ;
        RECT 9.100 0.530 12.625 0.760 ;
        RECT 16.595 0.740 16.825 1.435 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnrnq_4
MACRO gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.080 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.433000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.890 1.770 4.050 2.150 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.284000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.380 1.770 20.630 2.150 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.149500 ;
    PORT
      LAYER Metal1 ;
        RECT 17.450 1.770 18.550 2.150 ;
        RECT 18.280 1.320 18.550 1.770 ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.675500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.280 1.770 1.590 2.150 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.895400 ;
    PORT
      LAYER Metal1 ;
        RECT 23.585 0.550 23.960 3.380 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 24.080 4.220 ;
        RECT 1.310 3.005 1.650 3.620 ;
        RECT 3.050 3.000 3.390 3.620 ;
        RECT 7.585 3.165 7.930 3.620 ;
        RECT 13.450 3.035 13.680 3.620 ;
        RECT 17.705 2.940 18.045 3.620 ;
        RECT 19.745 2.940 20.085 3.620 ;
        RECT 21.840 2.415 22.070 3.620 ;
        RECT 22.580 2.565 22.810 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.980 24.510 4.350 ;
        RECT -0.430 1.760 9.885 1.980 ;
        RECT 17.020 1.760 24.510 1.980 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 9.885 1.760 17.020 1.980 ;
        RECT -0.430 -0.430 24.510 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 1.050 ;
        RECT 3.270 0.300 3.610 1.075 ;
        RECT 10.580 0.300 10.920 0.915 ;
        RECT 19.745 0.300 20.085 1.075 ;
        RECT 22.480 0.300 22.710 0.930 ;
        RECT 0.000 -0.300 24.080 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 2.670 0.575 3.300 ;
        RECT 2.385 2.770 2.615 3.300 ;
        RECT 3.785 3.105 7.095 3.335 ;
        RECT 3.785 2.770 4.015 3.105 ;
        RECT 6.865 2.935 7.095 3.105 ;
        RECT 8.280 3.160 13.220 3.390 ;
        RECT 8.280 2.935 8.510 3.160 ;
        RECT 0.345 2.435 2.055 2.670 ;
        RECT 1.825 1.510 2.055 2.435 ;
        RECT 0.245 1.280 2.055 1.510 ;
        RECT 2.385 2.540 4.015 2.770 ;
        RECT 0.245 0.810 0.475 1.280 ;
        RECT 2.385 1.150 2.615 2.540 ;
        RECT 2.385 0.810 2.715 1.150 ;
        RECT 4.290 0.845 4.730 2.830 ;
        RECT 5.310 2.015 5.650 2.830 ;
        RECT 6.405 2.475 6.635 2.870 ;
        RECT 6.865 2.705 8.510 2.935 ;
        RECT 10.510 2.815 10.850 2.875 ;
        RECT 8.740 2.585 10.850 2.815 ;
        RECT 11.790 2.645 12.760 2.875 ;
        RECT 8.740 2.475 8.970 2.585 ;
        RECT 6.405 2.245 8.970 2.475 ;
        RECT 12.530 2.345 12.760 2.645 ;
        RECT 12.990 2.805 13.220 3.160 ;
        RECT 14.175 3.160 15.480 3.390 ;
        RECT 14.175 2.805 14.405 3.160 ;
        RECT 12.990 2.575 14.405 2.805 ;
        RECT 14.635 2.345 14.975 2.875 ;
        RECT 9.200 2.070 12.300 2.300 ;
        RECT 12.530 2.125 14.975 2.345 ;
        RECT 12.530 2.115 14.750 2.125 ;
        RECT 9.200 2.015 9.430 2.070 ;
        RECT 5.310 1.785 9.430 2.015 ;
        RECT 5.565 0.790 5.795 1.785 ;
        RECT 9.660 1.605 11.840 1.835 ;
        RECT 9.660 1.555 9.890 1.605 ;
        RECT 6.135 1.020 6.475 1.555 ;
        RECT 7.030 1.325 9.890 1.555 ;
        RECT 10.120 1.145 11.380 1.375 ;
        RECT 10.120 1.020 10.350 1.145 ;
        RECT 6.135 0.790 10.350 1.020 ;
        RECT 11.150 0.760 11.380 1.145 ;
        RECT 11.610 1.315 11.840 1.605 ;
        RECT 12.070 1.775 12.300 2.070 ;
        RECT 12.070 1.545 12.470 1.775 ;
        RECT 14.465 1.315 14.750 2.115 ;
        RECT 15.250 2.070 15.480 3.160 ;
        RECT 15.710 3.160 17.475 3.390 ;
        RECT 15.710 1.315 15.940 3.160 ;
        RECT 16.675 1.370 17.015 2.895 ;
        RECT 17.245 2.710 17.475 3.160 ;
        RECT 18.275 3.085 19.470 3.320 ;
        RECT 18.275 2.710 18.505 3.085 ;
        RECT 17.245 2.475 18.505 2.710 ;
        RECT 11.610 1.085 14.750 1.315 ;
        RECT 14.980 1.085 15.940 1.315 ;
        RECT 16.170 1.315 17.015 1.370 ;
        RECT 16.170 1.085 17.925 1.315 ;
        RECT 16.170 1.030 16.455 1.085 ;
        RECT 17.640 1.075 17.925 1.085 ;
        RECT 18.780 1.075 19.010 2.855 ;
        RECT 19.240 2.710 19.470 3.085 ;
        RECT 20.315 3.085 21.610 3.320 ;
        RECT 20.315 2.710 20.545 3.085 ;
        RECT 19.240 2.480 20.545 2.710 ;
        RECT 20.820 2.515 21.150 2.855 ;
        RECT 20.920 1.560 21.150 2.515 ;
        RECT 21.380 1.910 21.610 3.085 ;
        RECT 20.920 1.540 23.250 1.560 ;
        RECT 19.305 1.330 23.250 1.540 ;
        RECT 19.305 1.310 21.990 1.330 ;
        RECT 14.430 0.760 14.770 0.855 ;
        RECT 16.775 0.760 17.115 0.855 ;
        RECT 17.640 0.790 19.010 1.075 ;
        RECT 21.760 0.790 21.990 1.310 ;
        RECT 11.150 0.530 17.115 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_1
MACRO gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.200 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.433000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.890 1.770 4.050 2.150 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.284000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.380 1.770 20.630 2.150 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.149500 ;
    PORT
      LAYER Metal1 ;
        RECT 17.450 1.770 18.540 2.150 ;
        RECT 18.225 1.340 18.540 1.770 ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.675500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.280 1.770 1.590 2.150 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.058200 ;
    PORT
      LAYER Metal1 ;
        RECT 23.545 2.320 23.980 3.380 ;
        RECT 23.545 2.070 24.550 2.320 ;
        RECT 24.170 1.170 24.550 2.070 ;
        RECT 23.600 0.940 24.550 1.170 ;
        RECT 23.600 0.550 23.980 0.940 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 25.200 4.220 ;
        RECT 1.310 3.005 1.650 3.620 ;
        RECT 3.050 3.000 3.390 3.620 ;
        RECT 7.585 3.165 7.930 3.620 ;
        RECT 13.450 3.035 13.680 3.620 ;
        RECT 17.705 2.940 18.045 3.620 ;
        RECT 19.745 2.940 20.085 3.620 ;
        RECT 21.840 2.415 22.070 3.620 ;
        RECT 22.580 2.570 22.810 3.620 ;
        RECT 24.620 2.570 24.850 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.980 25.630 4.350 ;
        RECT -0.430 1.760 9.885 1.980 ;
        RECT 17.020 1.760 25.630 1.980 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 9.885 1.760 17.020 1.980 ;
        RECT -0.430 -0.430 25.630 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 1.050 ;
        RECT 3.270 0.300 3.610 1.075 ;
        RECT 10.580 0.300 10.920 0.915 ;
        RECT 19.745 0.300 20.085 1.075 ;
        RECT 22.480 0.300 22.710 0.765 ;
        RECT 24.665 0.300 25.005 0.710 ;
        RECT 0.000 -0.300 25.200 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 2.670 0.575 3.300 ;
        RECT 2.385 2.770 2.615 3.300 ;
        RECT 3.785 3.105 7.095 3.335 ;
        RECT 3.785 2.770 4.015 3.105 ;
        RECT 6.865 2.935 7.095 3.105 ;
        RECT 8.280 3.160 13.220 3.390 ;
        RECT 8.280 2.935 8.510 3.160 ;
        RECT 0.345 2.435 2.055 2.670 ;
        RECT 1.825 1.510 2.055 2.435 ;
        RECT 0.245 1.280 2.055 1.510 ;
        RECT 2.385 2.540 4.015 2.770 ;
        RECT 0.245 0.810 0.475 1.280 ;
        RECT 2.385 1.150 2.615 2.540 ;
        RECT 2.385 0.810 2.715 1.150 ;
        RECT 4.290 0.845 4.730 2.830 ;
        RECT 5.310 2.015 5.650 2.830 ;
        RECT 6.405 2.475 6.635 2.870 ;
        RECT 6.865 2.705 8.510 2.935 ;
        RECT 10.510 2.815 10.850 2.875 ;
        RECT 8.740 2.585 10.850 2.815 ;
        RECT 11.790 2.645 12.760 2.875 ;
        RECT 8.740 2.475 8.970 2.585 ;
        RECT 6.405 2.245 8.970 2.475 ;
        RECT 12.530 2.345 12.760 2.645 ;
        RECT 12.990 2.805 13.220 3.160 ;
        RECT 14.175 3.160 15.480 3.390 ;
        RECT 14.175 2.805 14.405 3.160 ;
        RECT 12.990 2.575 14.405 2.805 ;
        RECT 14.635 2.345 14.975 2.875 ;
        RECT 9.200 2.070 12.300 2.300 ;
        RECT 12.530 2.125 14.975 2.345 ;
        RECT 12.530 2.115 14.750 2.125 ;
        RECT 9.200 2.015 9.430 2.070 ;
        RECT 5.310 1.785 9.430 2.015 ;
        RECT 5.565 0.790 5.795 1.785 ;
        RECT 9.660 1.605 11.840 1.835 ;
        RECT 9.660 1.555 9.890 1.605 ;
        RECT 6.135 1.020 6.475 1.555 ;
        RECT 7.030 1.325 9.890 1.555 ;
        RECT 10.120 1.145 11.380 1.375 ;
        RECT 10.120 1.020 10.350 1.145 ;
        RECT 6.135 0.790 10.350 1.020 ;
        RECT 11.150 0.760 11.380 1.145 ;
        RECT 11.610 1.315 11.840 1.605 ;
        RECT 12.070 1.775 12.300 2.070 ;
        RECT 12.070 1.545 12.470 1.775 ;
        RECT 14.465 1.315 14.750 2.115 ;
        RECT 15.250 2.070 15.480 3.160 ;
        RECT 15.710 3.160 17.475 3.390 ;
        RECT 15.710 1.315 15.940 3.160 ;
        RECT 16.675 1.370 17.015 2.895 ;
        RECT 17.245 2.710 17.475 3.160 ;
        RECT 18.275 3.085 19.470 3.320 ;
        RECT 18.275 2.710 18.505 3.085 ;
        RECT 17.245 2.475 18.505 2.710 ;
        RECT 11.610 1.085 14.750 1.315 ;
        RECT 14.980 1.085 15.940 1.315 ;
        RECT 16.170 1.315 17.015 1.370 ;
        RECT 16.170 1.085 17.995 1.315 ;
        RECT 16.170 1.030 16.455 1.085 ;
        RECT 17.710 1.075 17.995 1.085 ;
        RECT 18.780 1.075 19.010 2.855 ;
        RECT 19.240 2.710 19.470 3.085 ;
        RECT 20.315 3.085 21.610 3.320 ;
        RECT 20.315 2.710 20.545 3.085 ;
        RECT 19.240 2.480 20.545 2.710 ;
        RECT 20.820 2.515 21.150 2.855 ;
        RECT 20.920 1.560 21.150 2.515 ;
        RECT 21.380 1.910 21.610 3.085 ;
        RECT 22.965 1.560 23.720 1.820 ;
        RECT 20.920 1.540 23.720 1.560 ;
        RECT 19.305 1.475 23.720 1.540 ;
        RECT 19.305 1.330 23.305 1.475 ;
        RECT 19.305 1.310 21.990 1.330 ;
        RECT 14.430 0.760 14.770 0.855 ;
        RECT 16.775 0.760 17.115 0.855 ;
        RECT 17.710 0.790 19.010 1.075 ;
        RECT 21.760 0.790 21.990 1.310 ;
        RECT 11.150 0.530 17.115 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_2
MACRO gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.440 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.433000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.890 1.770 4.050 2.150 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.284000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.380 1.770 20.630 2.150 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.149500 ;
    PORT
      LAYER Metal1 ;
        RECT 17.450 1.770 18.540 2.150 ;
        RECT 18.225 1.320 18.540 1.770 ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.675500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.280 1.770 1.590 2.150 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.111200 ;
    PORT
      LAYER Metal1 ;
        RECT 23.545 2.330 23.885 3.380 ;
        RECT 25.585 2.330 26.230 3.380 ;
        RECT 23.545 2.100 26.230 2.330 ;
        RECT 25.850 1.170 26.230 2.100 ;
        RECT 23.600 0.940 26.230 1.170 ;
        RECT 23.600 0.550 23.830 0.940 ;
        RECT 25.840 0.550 26.230 0.940 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 27.440 4.220 ;
        RECT 1.310 3.005 1.650 3.620 ;
        RECT 3.050 3.000 3.390 3.620 ;
        RECT 7.585 3.165 7.930 3.620 ;
        RECT 13.450 3.035 13.680 3.620 ;
        RECT 17.705 2.940 18.045 3.620 ;
        RECT 19.745 2.940 20.085 3.620 ;
        RECT 21.840 2.415 22.070 3.620 ;
        RECT 22.580 2.570 22.810 3.620 ;
        RECT 24.620 2.570 24.850 3.620 ;
        RECT 26.660 2.570 26.890 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.980 27.870 4.350 ;
        RECT -0.430 1.760 9.885 1.980 ;
        RECT 17.020 1.760 27.870 1.980 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 9.885 1.760 17.020 1.980 ;
        RECT -0.430 -0.430 27.870 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 1.050 ;
        RECT 3.270 0.300 3.610 1.075 ;
        RECT 10.580 0.300 10.920 0.915 ;
        RECT 19.745 0.300 20.085 1.075 ;
        RECT 22.480 0.300 22.710 0.765 ;
        RECT 24.665 0.300 25.005 0.710 ;
        RECT 26.960 0.300 27.190 0.765 ;
        RECT 0.000 -0.300 27.440 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 2.670 0.575 3.300 ;
        RECT 2.385 2.770 2.615 3.300 ;
        RECT 3.785 3.105 7.095 3.335 ;
        RECT 3.785 2.770 4.015 3.105 ;
        RECT 6.865 2.935 7.095 3.105 ;
        RECT 8.280 3.160 13.220 3.390 ;
        RECT 8.280 2.935 8.510 3.160 ;
        RECT 0.345 2.435 2.055 2.670 ;
        RECT 1.825 1.510 2.055 2.435 ;
        RECT 0.245 1.280 2.055 1.510 ;
        RECT 2.385 2.540 4.015 2.770 ;
        RECT 0.245 0.810 0.475 1.280 ;
        RECT 2.385 1.150 2.615 2.540 ;
        RECT 2.385 0.810 2.715 1.150 ;
        RECT 4.290 0.845 4.730 2.830 ;
        RECT 5.310 2.015 5.650 2.830 ;
        RECT 6.405 2.475 6.635 2.870 ;
        RECT 6.865 2.705 8.510 2.935 ;
        RECT 10.510 2.815 10.850 2.875 ;
        RECT 8.740 2.585 10.850 2.815 ;
        RECT 11.790 2.645 12.760 2.875 ;
        RECT 8.740 2.475 8.970 2.585 ;
        RECT 6.405 2.245 8.970 2.475 ;
        RECT 12.530 2.345 12.760 2.645 ;
        RECT 12.990 2.805 13.220 3.160 ;
        RECT 14.175 3.160 15.480 3.390 ;
        RECT 14.175 2.805 14.405 3.160 ;
        RECT 12.990 2.575 14.405 2.805 ;
        RECT 14.635 2.345 14.975 2.875 ;
        RECT 9.200 2.070 12.300 2.300 ;
        RECT 12.530 2.125 14.975 2.345 ;
        RECT 12.530 2.115 14.750 2.125 ;
        RECT 9.200 2.015 9.430 2.070 ;
        RECT 5.310 1.785 9.430 2.015 ;
        RECT 5.565 0.790 5.795 1.785 ;
        RECT 9.660 1.605 11.840 1.835 ;
        RECT 9.660 1.555 9.890 1.605 ;
        RECT 6.135 1.020 6.475 1.555 ;
        RECT 7.030 1.325 9.890 1.555 ;
        RECT 10.120 1.145 11.380 1.375 ;
        RECT 10.120 1.020 10.350 1.145 ;
        RECT 6.135 0.790 10.350 1.020 ;
        RECT 11.150 0.760 11.380 1.145 ;
        RECT 11.610 1.315 11.840 1.605 ;
        RECT 12.070 1.775 12.300 2.070 ;
        RECT 12.070 1.545 12.470 1.775 ;
        RECT 14.465 1.315 14.750 2.115 ;
        RECT 15.250 2.070 15.480 3.160 ;
        RECT 15.710 3.160 17.475 3.390 ;
        RECT 15.710 1.315 15.940 3.160 ;
        RECT 16.675 1.370 17.015 2.895 ;
        RECT 17.245 2.710 17.475 3.160 ;
        RECT 18.275 3.085 19.470 3.320 ;
        RECT 18.275 2.710 18.505 3.085 ;
        RECT 17.245 2.475 18.505 2.710 ;
        RECT 11.610 1.085 14.750 1.315 ;
        RECT 14.980 1.085 15.940 1.315 ;
        RECT 16.170 1.315 17.015 1.370 ;
        RECT 16.170 1.085 17.960 1.315 ;
        RECT 16.170 1.030 16.455 1.085 ;
        RECT 17.675 1.075 17.960 1.085 ;
        RECT 18.780 1.075 19.010 2.855 ;
        RECT 19.240 2.710 19.470 3.085 ;
        RECT 20.315 3.085 21.610 3.320 ;
        RECT 20.315 2.710 20.545 3.085 ;
        RECT 19.240 2.480 20.545 2.710 ;
        RECT 20.820 2.515 21.150 2.855 ;
        RECT 20.920 1.560 21.150 2.515 ;
        RECT 21.380 1.910 21.610 3.085 ;
        RECT 22.965 1.560 25.390 1.820 ;
        RECT 20.920 1.540 25.390 1.560 ;
        RECT 19.305 1.475 25.390 1.540 ;
        RECT 19.305 1.330 23.305 1.475 ;
        RECT 19.305 1.310 21.990 1.330 ;
        RECT 14.430 0.760 14.770 0.855 ;
        RECT 16.775 0.760 17.115 0.855 ;
        RECT 17.675 0.790 19.010 1.075 ;
        RECT 21.760 0.790 21.990 1.310 ;
        RECT 11.150 0.530 17.115 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_4
MACRO gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.160 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.530500 ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 1.770 4.390 2.150 ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.156500 ;
    PORT
      LAYER Metal1 ;
        RECT 14.560 1.220 15.590 1.670 ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.794000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.280 1.770 1.590 2.130 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.893200 ;
    PORT
      LAYER Metal1 ;
        RECT 19.610 0.550 20.040 3.380 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 20.160 4.220 ;
        RECT 1.310 3.005 1.650 3.620 ;
        RECT 3.050 3.005 3.390 3.620 ;
        RECT 7.290 3.240 7.630 3.620 ;
        RECT 9.825 2.885 10.055 3.620 ;
        RECT 14.110 2.945 14.450 3.620 ;
        RECT 16.745 2.600 16.975 3.620 ;
        RECT 18.645 2.530 18.875 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 20.590 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 20.590 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.935 ;
        RECT 3.225 0.300 3.455 1.145 ;
        RECT 7.470 0.300 7.810 1.090 ;
        RECT 16.650 0.300 16.990 1.080 ;
        RECT 18.545 0.300 18.775 0.835 ;
        RECT 0.000 -0.300 20.160 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 2.595 0.575 3.300 ;
        RECT 2.385 2.775 2.715 3.300 ;
        RECT 3.620 3.120 6.230 3.360 ;
        RECT 3.620 2.775 3.850 3.120 ;
        RECT 0.345 2.360 2.155 2.595 ;
        RECT 1.925 1.395 2.155 2.360 ;
        RECT 0.245 1.165 2.155 1.395 ;
        RECT 2.385 2.545 3.850 2.775 ;
        RECT 5.940 2.880 6.230 3.120 ;
        RECT 7.975 2.885 9.330 3.115 ;
        RECT 7.975 2.880 8.205 2.885 ;
        RECT 0.245 0.660 0.475 1.165 ;
        RECT 2.385 0.660 2.715 2.545 ;
        RECT 4.290 2.520 5.090 2.750 ;
        RECT 4.860 1.095 5.090 2.520 ;
        RECT 4.290 0.865 5.090 1.095 ;
        RECT 5.365 1.630 5.595 2.710 ;
        RECT 5.940 2.650 8.205 2.880 ;
        RECT 9.100 2.655 9.330 2.885 ;
        RECT 10.285 3.065 11.670 3.295 ;
        RECT 10.285 2.655 10.515 3.065 ;
        RECT 12.145 2.940 13.855 3.175 ;
        RECT 8.530 2.195 8.870 2.655 ;
        RECT 9.100 2.425 10.515 2.655 ;
        RECT 10.890 2.195 11.230 2.655 ;
        RECT 6.630 1.965 11.230 2.195 ;
        RECT 9.825 1.930 11.230 1.965 ;
        RECT 5.365 1.395 8.290 1.630 ;
        RECT 5.365 0.865 5.850 1.395 ;
        RECT 9.825 0.810 10.055 1.930 ;
        RECT 12.145 1.585 12.375 2.940 ;
        RECT 13.625 2.715 13.855 2.940 ;
        RECT 14.755 2.885 16.380 3.120 ;
        RECT 14.755 2.715 14.985 2.885 ;
        RECT 10.945 1.355 12.375 1.585 ;
        RECT 13.165 2.195 13.395 2.710 ;
        RECT 13.625 2.480 14.985 2.715 ;
        RECT 15.380 2.195 15.730 2.655 ;
        RECT 13.165 1.965 15.730 2.195 ;
        RECT 16.150 2.195 16.380 2.885 ;
        RECT 10.945 0.810 11.175 1.355 ;
        RECT 13.165 1.135 13.395 1.965 ;
        RECT 16.150 1.960 17.470 2.195 ;
        RECT 17.765 1.895 17.995 2.875 ;
        RECT 17.765 1.615 19.215 1.895 ;
        RECT 15.990 1.545 19.215 1.615 ;
        RECT 15.990 1.385 18.055 1.545 ;
        RECT 13.165 1.075 14.295 1.135 ;
        RECT 12.010 0.795 14.295 1.075 ;
        RECT 17.825 0.795 18.055 1.385 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1
MACRO gf180mcu_fd_sc_mcu7t5v0__dffnsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.530500 ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 1.770 4.390 2.150 ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.156500 ;
    PORT
      LAYER Metal1 ;
        RECT 14.560 1.220 15.590 1.670 ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.794000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.280 1.770 1.590 2.130 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.055600 ;
    PORT
      LAYER Metal1 ;
        RECT 19.610 2.320 20.060 3.380 ;
        RECT 19.610 2.090 20.620 2.320 ;
        RECT 20.260 1.290 20.620 2.090 ;
        RECT 19.665 1.060 20.620 1.290 ;
        RECT 19.665 0.550 20.060 1.060 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 21.280 4.220 ;
        RECT 1.310 3.005 1.650 3.620 ;
        RECT 3.050 3.005 3.390 3.620 ;
        RECT 7.290 3.240 7.630 3.620 ;
        RECT 9.825 2.885 10.055 3.620 ;
        RECT 14.110 2.945 14.450 3.620 ;
        RECT 16.745 2.600 16.975 3.620 ;
        RECT 18.645 2.570 18.875 3.620 ;
        RECT 20.685 2.570 20.915 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 21.710 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.710 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.935 ;
        RECT 3.225 0.300 3.455 1.145 ;
        RECT 7.470 0.300 7.810 1.090 ;
        RECT 16.650 0.300 16.990 1.080 ;
        RECT 18.545 0.300 18.775 0.765 ;
        RECT 20.785 0.300 21.015 0.765 ;
        RECT 0.000 -0.300 21.280 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 2.595 0.575 3.300 ;
        RECT 2.385 2.775 2.715 3.300 ;
        RECT 3.620 3.120 6.230 3.360 ;
        RECT 3.620 2.775 3.850 3.120 ;
        RECT 0.345 2.360 2.155 2.595 ;
        RECT 1.925 1.395 2.155 2.360 ;
        RECT 0.245 1.165 2.155 1.395 ;
        RECT 2.385 2.545 3.850 2.775 ;
        RECT 5.940 2.880 6.230 3.120 ;
        RECT 7.975 2.885 9.330 3.115 ;
        RECT 7.975 2.880 8.205 2.885 ;
        RECT 0.245 0.660 0.475 1.165 ;
        RECT 2.385 0.660 2.715 2.545 ;
        RECT 4.290 2.520 5.090 2.750 ;
        RECT 4.860 1.095 5.090 2.520 ;
        RECT 4.290 0.865 5.090 1.095 ;
        RECT 5.365 1.630 5.595 2.710 ;
        RECT 5.940 2.650 8.205 2.880 ;
        RECT 9.100 2.655 9.330 2.885 ;
        RECT 10.285 3.065 11.670 3.295 ;
        RECT 10.285 2.655 10.515 3.065 ;
        RECT 12.145 2.940 13.855 3.175 ;
        RECT 8.530 2.195 8.870 2.655 ;
        RECT 9.100 2.425 10.515 2.655 ;
        RECT 10.890 2.195 11.230 2.655 ;
        RECT 6.630 1.965 11.230 2.195 ;
        RECT 9.825 1.930 11.230 1.965 ;
        RECT 5.365 1.395 8.290 1.630 ;
        RECT 5.365 0.865 5.850 1.395 ;
        RECT 9.825 0.810 10.055 1.930 ;
        RECT 12.145 1.585 12.375 2.940 ;
        RECT 13.625 2.715 13.855 2.940 ;
        RECT 14.755 2.885 16.380 3.120 ;
        RECT 14.755 2.715 14.985 2.885 ;
        RECT 10.945 1.355 12.375 1.585 ;
        RECT 13.165 2.195 13.395 2.710 ;
        RECT 13.625 2.480 14.985 2.715 ;
        RECT 15.380 2.195 15.730 2.655 ;
        RECT 13.165 1.965 15.730 2.195 ;
        RECT 16.150 2.195 16.380 2.885 ;
        RECT 10.945 0.810 11.175 1.355 ;
        RECT 13.165 1.135 13.395 1.965 ;
        RECT 16.150 1.960 17.470 2.195 ;
        RECT 17.765 1.835 17.995 2.875 ;
        RECT 17.765 1.615 19.930 1.835 ;
        RECT 15.990 1.605 19.930 1.615 ;
        RECT 15.990 1.385 18.055 1.605 ;
        RECT 13.165 1.075 14.295 1.135 ;
        RECT 12.010 0.795 14.295 1.075 ;
        RECT 17.825 0.795 18.055 1.385 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnsnq_2
MACRO gf180mcu_fd_sc_mcu7t5v0__dffnsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.520 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.530500 ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 1.770 4.390 2.150 ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.156500 ;
    PORT
      LAYER Metal1 ;
        RECT 14.560 1.220 15.590 1.670 ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.794000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.280 1.770 1.590 2.130 ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.111200 ;
    PORT
      LAYER Metal1 ;
        RECT 19.665 2.320 19.895 3.380 ;
        RECT 21.690 2.320 22.310 3.380 ;
        RECT 19.665 2.090 22.310 2.320 ;
        RECT 21.930 1.290 22.310 2.090 ;
        RECT 19.665 1.060 22.310 1.290 ;
        RECT 19.665 0.805 19.895 1.060 ;
        RECT 21.905 0.550 22.310 1.060 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 23.520 4.220 ;
        RECT 1.310 3.005 1.650 3.620 ;
        RECT 3.050 3.005 3.390 3.620 ;
        RECT 7.290 3.240 7.630 3.620 ;
        RECT 9.825 2.885 10.055 3.620 ;
        RECT 14.110 2.945 14.450 3.620 ;
        RECT 16.745 2.600 16.975 3.620 ;
        RECT 18.645 2.570 18.875 3.620 ;
        RECT 20.685 2.570 20.915 3.620 ;
        RECT 22.725 2.570 22.955 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 23.950 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 23.950 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.935 ;
        RECT 3.225 0.300 3.455 1.145 ;
        RECT 7.470 0.300 7.810 1.090 ;
        RECT 16.650 0.300 16.990 1.080 ;
        RECT 18.545 0.300 18.775 0.765 ;
        RECT 20.785 0.300 21.015 0.765 ;
        RECT 23.025 0.300 23.255 0.765 ;
        RECT 0.000 -0.300 23.520 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 2.595 0.575 3.300 ;
        RECT 2.385 2.775 2.715 3.300 ;
        RECT 3.620 3.120 6.230 3.360 ;
        RECT 3.620 2.775 3.850 3.120 ;
        RECT 0.345 2.360 2.155 2.595 ;
        RECT 1.925 1.395 2.155 2.360 ;
        RECT 0.245 1.165 2.155 1.395 ;
        RECT 2.385 2.545 3.850 2.775 ;
        RECT 5.940 2.880 6.230 3.120 ;
        RECT 7.975 2.885 9.330 3.115 ;
        RECT 7.975 2.880 8.205 2.885 ;
        RECT 0.245 0.660 0.475 1.165 ;
        RECT 2.385 0.660 2.715 2.545 ;
        RECT 4.290 2.520 5.090 2.750 ;
        RECT 4.860 1.095 5.090 2.520 ;
        RECT 4.290 0.865 5.090 1.095 ;
        RECT 5.365 1.630 5.595 2.710 ;
        RECT 5.940 2.650 8.205 2.880 ;
        RECT 9.100 2.655 9.330 2.885 ;
        RECT 10.285 3.065 11.670 3.295 ;
        RECT 10.285 2.655 10.515 3.065 ;
        RECT 12.145 2.940 13.855 3.175 ;
        RECT 8.530 2.195 8.870 2.655 ;
        RECT 9.100 2.425 10.515 2.655 ;
        RECT 10.890 2.195 11.230 2.655 ;
        RECT 6.630 1.965 11.230 2.195 ;
        RECT 9.825 1.930 11.230 1.965 ;
        RECT 5.365 1.395 8.290 1.630 ;
        RECT 5.365 0.865 5.850 1.395 ;
        RECT 9.825 0.810 10.055 1.930 ;
        RECT 12.145 1.585 12.375 2.940 ;
        RECT 13.625 2.715 13.855 2.940 ;
        RECT 14.755 2.885 16.380 3.120 ;
        RECT 14.755 2.715 14.985 2.885 ;
        RECT 10.945 1.355 12.375 1.585 ;
        RECT 13.165 2.195 13.395 2.710 ;
        RECT 13.625 2.480 14.985 2.715 ;
        RECT 15.380 2.195 15.730 2.655 ;
        RECT 13.165 1.965 15.730 2.195 ;
        RECT 16.150 2.195 16.380 2.885 ;
        RECT 10.945 0.810 11.175 1.355 ;
        RECT 13.165 1.135 13.395 1.965 ;
        RECT 16.150 1.960 17.470 2.195 ;
        RECT 17.765 1.840 17.995 2.875 ;
        RECT 17.765 1.615 21.560 1.840 ;
        RECT 15.990 1.605 21.560 1.615 ;
        RECT 15.990 1.385 18.055 1.605 ;
        RECT 13.165 1.075 14.295 1.135 ;
        RECT 12.010 0.795 14.295 1.075 ;
        RECT 17.825 0.795 18.055 1.385 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnsnq_4
MACRO gf180mcu_fd_sc_mcu7t5v0__dffq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.240 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.570 1.210 4.975 2.710 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.675500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 1.770 1.590 2.150 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 14.835 2.330 15.850 2.975 ;
        RECT 15.470 0.550 15.850 2.330 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 16.240 4.220 ;
        RECT 1.310 2.930 1.650 3.620 ;
        RECT 3.305 3.185 3.535 3.620 ;
        RECT 7.630 2.700 7.970 3.620 ;
        RECT 12.625 2.635 12.855 3.620 ;
        RECT 14.365 2.635 14.595 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 16.670 4.350 ;
        RECT -0.430 1.760 4.865 1.885 ;
        RECT 6.120 1.760 16.670 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 4.865 1.760 6.120 1.885 ;
        RECT -0.430 -0.430 16.670 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 1.050 ;
        RECT 3.150 0.300 3.490 1.090 ;
        RECT 7.790 0.300 8.130 0.585 ;
        RECT 12.485 0.300 12.715 1.105 ;
        RECT 14.425 0.300 14.655 0.890 ;
        RECT 0.000 -0.300 16.240 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 2.700 0.575 3.155 ;
        RECT 1.915 2.980 3.075 3.215 ;
        RECT 1.915 2.700 2.145 2.980 ;
        RECT 2.845 2.885 3.075 2.980 ;
        RECT 3.890 3.160 6.590 3.390 ;
        RECT 8.640 3.160 11.330 3.390 ;
        RECT 3.890 2.885 4.120 3.160 ;
        RECT 0.345 2.470 2.145 2.700 ;
        RECT 1.915 1.510 2.145 2.470 ;
        RECT 2.385 2.325 2.615 2.710 ;
        RECT 2.845 2.650 4.120 2.885 ;
        RECT 5.610 2.470 5.950 2.930 ;
        RECT 2.385 2.090 4.075 2.325 ;
        RECT 3.845 1.555 4.075 2.090 ;
        RECT 0.245 1.280 2.145 1.510 ;
        RECT 2.485 1.325 4.075 1.555 ;
        RECT 0.245 0.810 0.475 1.280 ;
        RECT 2.485 0.810 2.715 1.325 ;
        RECT 3.845 0.760 4.075 1.325 ;
        RECT 5.325 2.240 8.410 2.470 ;
        RECT 5.325 0.990 5.670 2.240 ;
        RECT 8.640 2.010 8.870 3.160 ;
        RECT 6.165 1.780 8.870 2.010 ;
        RECT 6.165 0.760 6.395 1.780 ;
        RECT 9.125 1.550 9.470 2.930 ;
        RECT 7.130 1.320 9.470 1.550 ;
        RECT 9.130 0.860 9.470 1.320 ;
        RECT 9.720 1.225 9.950 3.160 ;
        RECT 10.250 2.130 10.590 2.930 ;
        RECT 10.250 1.895 13.350 2.130 ;
        RECT 10.250 0.860 10.590 1.895 ;
        RECT 13.645 1.840 13.875 3.030 ;
        RECT 13.645 1.630 15.095 1.840 ;
        RECT 11.770 1.500 15.095 1.630 ;
        RECT 11.770 1.400 13.870 1.500 ;
        RECT 3.845 0.530 6.395 0.760 ;
        RECT 13.605 0.755 13.870 1.400 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffq_1
MACRO gf180mcu_fd_sc_mcu7t5v0__dffq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.360 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.570 1.210 4.975 2.710 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.675500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 1.770 1.590 2.150 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.060800 ;
    PORT
      LAYER Metal1 ;
        RECT 15.330 2.330 16.410 2.975 ;
        RECT 16.030 1.020 16.410 2.330 ;
        RECT 15.450 0.550 16.410 1.020 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 17.360 4.220 ;
        RECT 1.310 2.930 1.650 3.620 ;
        RECT 3.305 3.185 3.535 3.620 ;
        RECT 7.630 2.700 7.970 3.620 ;
        RECT 12.625 2.635 12.855 3.620 ;
        RECT 14.365 2.635 14.595 3.620 ;
        RECT 16.665 2.635 16.895 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 17.790 4.350 ;
        RECT -0.430 1.760 4.865 1.885 ;
        RECT 6.120 1.760 17.790 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 4.865 1.760 6.120 1.885 ;
        RECT -0.430 -0.430 17.790 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 1.050 ;
        RECT 3.150 0.300 3.490 1.090 ;
        RECT 7.790 0.300 8.130 0.585 ;
        RECT 12.485 0.300 12.715 1.105 ;
        RECT 14.425 0.300 14.655 0.890 ;
        RECT 16.665 0.300 16.895 0.970 ;
        RECT 0.000 -0.300 17.360 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 2.700 0.575 3.155 ;
        RECT 1.915 2.980 3.075 3.215 ;
        RECT 1.915 2.700 2.145 2.980 ;
        RECT 2.845 2.885 3.075 2.980 ;
        RECT 3.890 3.160 6.590 3.390 ;
        RECT 8.640 3.160 11.330 3.390 ;
        RECT 3.890 2.885 4.120 3.160 ;
        RECT 0.345 2.470 2.145 2.700 ;
        RECT 1.915 1.510 2.145 2.470 ;
        RECT 2.385 2.325 2.615 2.710 ;
        RECT 2.845 2.650 4.120 2.885 ;
        RECT 5.610 2.470 5.950 2.930 ;
        RECT 2.385 2.090 4.075 2.325 ;
        RECT 3.845 1.555 4.075 2.090 ;
        RECT 0.245 1.280 2.145 1.510 ;
        RECT 2.485 1.325 4.075 1.555 ;
        RECT 0.245 0.810 0.475 1.280 ;
        RECT 2.485 0.810 2.715 1.325 ;
        RECT 3.845 0.760 4.075 1.325 ;
        RECT 5.325 2.240 8.410 2.470 ;
        RECT 5.325 0.990 5.670 2.240 ;
        RECT 8.640 2.010 8.870 3.160 ;
        RECT 6.165 1.780 8.870 2.010 ;
        RECT 6.165 0.760 6.395 1.780 ;
        RECT 9.125 1.550 9.470 2.930 ;
        RECT 7.130 1.320 9.470 1.550 ;
        RECT 9.130 0.860 9.470 1.320 ;
        RECT 9.720 1.225 9.950 3.160 ;
        RECT 10.250 2.130 10.590 2.930 ;
        RECT 10.250 1.895 13.350 2.130 ;
        RECT 10.250 0.860 10.590 1.895 ;
        RECT 13.645 1.840 13.875 3.030 ;
        RECT 13.645 1.630 15.565 1.840 ;
        RECT 11.770 1.500 15.565 1.630 ;
        RECT 11.770 1.400 13.870 1.500 ;
        RECT 13.605 0.805 13.870 1.400 ;
        RECT 3.845 0.530 6.395 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffq_2
MACRO gf180mcu_fd_sc_mcu7t5v0__dffq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.160 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.570 1.210 4.975 2.710 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.675500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.280 1.770 1.590 2.130 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.604400 ;
    PORT
      LAYER Metal1 ;
        RECT 15.735 2.330 18.510 2.930 ;
        RECT 18.130 1.170 18.510 2.330 ;
        RECT 15.965 0.940 18.510 1.170 ;
        RECT 15.965 0.805 16.195 0.940 ;
        RECT 17.795 0.835 18.510 0.940 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 20.160 4.220 ;
        RECT 1.310 2.930 1.650 3.620 ;
        RECT 3.305 3.185 3.535 3.620 ;
        RECT 7.630 2.700 7.970 3.620 ;
        RECT 12.625 2.720 12.855 3.620 ;
        RECT 14.725 2.720 14.955 3.620 ;
        RECT 17.030 3.285 17.370 3.620 ;
        RECT 19.325 2.720 19.555 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 20.590 4.350 ;
        RECT -0.430 1.760 4.865 1.885 ;
        RECT 6.120 1.760 20.590 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 4.865 1.760 6.120 1.885 ;
        RECT -0.430 -0.430 20.590 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 1.050 ;
        RECT 3.150 0.300 3.490 1.090 ;
        RECT 7.790 0.300 8.130 0.585 ;
        RECT 12.485 0.300 12.715 0.765 ;
        RECT 14.725 0.300 14.955 0.765 ;
        RECT 17.030 0.300 17.370 0.710 ;
        RECT 19.325 0.300 19.555 0.765 ;
        RECT 0.000 -0.300 20.160 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 2.590 0.575 3.225 ;
        RECT 1.915 2.980 3.075 3.215 ;
        RECT 1.915 2.590 2.145 2.980 ;
        RECT 2.845 2.885 3.075 2.980 ;
        RECT 3.890 3.160 6.590 3.390 ;
        RECT 8.640 3.160 11.330 3.390 ;
        RECT 3.890 2.885 4.120 3.160 ;
        RECT 0.345 2.360 2.145 2.590 ;
        RECT 1.915 1.510 2.145 2.360 ;
        RECT 2.385 2.325 2.615 2.710 ;
        RECT 2.845 2.650 4.120 2.885 ;
        RECT 5.610 2.470 5.950 2.930 ;
        RECT 2.385 2.090 4.075 2.325 ;
        RECT 3.845 1.555 4.075 2.090 ;
        RECT 0.245 1.280 2.145 1.510 ;
        RECT 2.485 1.325 4.075 1.555 ;
        RECT 0.245 0.810 0.475 1.280 ;
        RECT 2.485 0.810 2.715 1.325 ;
        RECT 3.845 0.760 4.075 1.325 ;
        RECT 5.325 2.240 8.410 2.470 ;
        RECT 5.325 0.990 5.670 2.240 ;
        RECT 8.640 2.010 8.870 3.160 ;
        RECT 6.165 1.780 8.870 2.010 ;
        RECT 6.165 0.760 6.395 1.780 ;
        RECT 9.125 1.550 9.470 2.930 ;
        RECT 7.130 1.320 9.470 1.550 ;
        RECT 9.130 0.860 9.470 1.320 ;
        RECT 9.720 1.225 9.950 3.160 ;
        RECT 10.250 2.130 10.590 2.930 ;
        RECT 10.250 1.895 13.350 2.130 ;
        RECT 10.250 0.860 10.590 1.895 ;
        RECT 13.645 1.840 13.875 3.070 ;
        RECT 13.645 1.630 17.795 1.840 ;
        RECT 11.770 1.500 17.795 1.630 ;
        RECT 11.770 1.400 13.870 1.500 ;
        RECT 13.605 0.805 13.870 1.400 ;
        RECT 3.845 0.530 6.395 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffq_4
MACRO gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.040 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.606000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.890 1.770 3.920 2.150 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.322000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.660 1.020 15.205 1.830 ;
        RECT 14.660 0.660 16.295 1.020 ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.675500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.280 1.770 1.570 2.150 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.893200 ;
    PORT
      LAYER Metal1 ;
        RECT 18.475 0.550 18.910 3.380 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 19.040 4.220 ;
        RECT 1.310 2.865 1.650 3.620 ;
        RECT 3.050 2.845 3.390 3.620 ;
        RECT 7.350 2.990 7.690 3.620 ;
        RECT 9.485 2.790 9.715 3.620 ;
        RECT 14.655 3.280 14.995 3.620 ;
        RECT 16.750 2.590 16.980 3.620 ;
        RECT 17.470 2.530 17.700 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.895 19.470 4.350 ;
        RECT -0.430 1.760 9.600 1.895 ;
        RECT 12.515 1.760 19.470 1.895 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 9.600 1.760 12.515 1.895 ;
        RECT -0.430 -0.430 19.470 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.655 1.050 ;
        RECT 3.170 0.300 3.510 1.075 ;
        RECT 8.430 0.300 8.770 0.915 ;
        RECT 14.070 0.300 14.300 1.130 ;
        RECT 17.315 0.300 17.655 0.875 ;
        RECT 0.000 -0.300 19.040 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 2.635 0.575 3.225 ;
        RECT 0.345 2.405 2.035 2.635 ;
        RECT 1.805 1.510 2.035 2.405 ;
        RECT 0.245 1.280 2.035 1.510 ;
        RECT 2.265 2.615 2.615 3.215 ;
        RECT 3.665 2.990 4.915 3.220 ;
        RECT 12.210 3.160 14.425 3.390 ;
        RECT 3.665 2.615 3.895 2.990 ;
        RECT 2.265 2.385 3.895 2.615 ;
        RECT 4.125 2.420 4.455 2.760 ;
        RECT 0.245 0.810 0.475 1.280 ;
        RECT 2.265 1.095 2.495 2.385 ;
        RECT 2.265 0.865 2.770 1.095 ;
        RECT 4.225 1.075 4.455 2.420 ;
        RECT 4.685 1.910 4.915 2.990 ;
        RECT 6.165 2.760 6.395 2.955 ;
        RECT 8.765 2.760 8.995 3.130 ;
        RECT 5.145 2.300 5.375 2.760 ;
        RECT 6.165 2.530 8.995 2.760 ;
        RECT 10.440 2.845 11.080 3.075 ;
        RECT 9.855 2.300 10.155 2.525 ;
        RECT 5.145 2.070 10.155 2.300 ;
        RECT 4.225 0.845 4.630 1.075 ;
        RECT 5.465 0.790 5.695 2.070 ;
        RECT 10.440 1.840 10.670 2.845 ;
        RECT 12.210 2.050 12.440 3.160 ;
        RECT 14.195 3.050 14.425 3.160 ;
        RECT 15.235 3.160 16.420 3.390 ;
        RECT 15.235 3.050 15.465 3.160 ;
        RECT 6.690 1.610 10.670 1.840 ;
        RECT 11.550 1.820 12.440 2.050 ;
        RECT 6.045 1.380 6.275 1.590 ;
        RECT 6.045 1.150 9.230 1.380 ;
        RECT 9.000 0.760 9.230 1.150 ;
        RECT 9.990 1.000 10.330 1.610 ;
        RECT 10.925 0.760 11.155 1.590 ;
        RECT 11.550 1.000 11.890 1.820 ;
        RECT 12.890 1.590 13.120 2.525 ;
        RECT 12.120 1.360 13.120 1.590 ;
        RECT 12.120 0.760 12.350 1.360 ;
        RECT 13.415 1.130 13.755 2.930 ;
        RECT 14.195 2.820 15.465 3.050 ;
        RECT 15.730 2.405 15.960 2.930 ;
        RECT 13.995 2.175 15.960 2.405 ;
        RECT 15.730 1.680 15.960 2.175 ;
        RECT 16.190 1.910 16.420 3.160 ;
        RECT 15.730 1.450 18.230 1.680 ;
        RECT 12.950 0.790 13.755 1.130 ;
        RECT 16.650 0.790 16.880 1.450 ;
        RECT 9.000 0.530 12.350 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
MACRO gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.160 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.606000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.890 1.770 3.920 2.150 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.429500 ;
    PORT
      LAYER Metal1 ;
        RECT 14.660 1.020 15.205 1.830 ;
        RECT 14.660 0.660 16.255 1.020 ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.675500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.280 1.770 1.570 2.150 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.055600 ;
    PORT
      LAYER Metal1 ;
        RECT 18.475 2.280 18.940 3.380 ;
        RECT 18.475 2.050 19.500 2.280 ;
        RECT 19.140 1.270 19.500 2.050 ;
        RECT 18.475 1.040 19.500 1.270 ;
        RECT 18.475 0.550 18.940 1.040 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 20.160 4.220 ;
        RECT 1.310 2.865 1.650 3.620 ;
        RECT 3.050 2.845 3.390 3.620 ;
        RECT 7.350 2.990 7.690 3.620 ;
        RECT 9.485 2.790 9.715 3.620 ;
        RECT 14.655 3.280 14.995 3.620 ;
        RECT 16.750 2.570 16.985 3.620 ;
        RECT 17.465 2.570 17.700 3.620 ;
        RECT 19.455 2.530 19.795 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.895 20.590 4.350 ;
        RECT -0.430 1.760 9.600 1.895 ;
        RECT 12.515 1.760 20.590 1.895 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 9.600 1.760 12.515 1.895 ;
        RECT -0.430 -0.430 20.590 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.655 1.050 ;
        RECT 3.170 0.300 3.510 1.075 ;
        RECT 8.430 0.300 8.770 0.915 ;
        RECT 14.070 0.300 14.300 1.130 ;
        RECT 17.315 0.300 17.655 0.790 ;
        RECT 19.555 0.300 19.895 0.790 ;
        RECT 0.000 -0.300 20.160 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 2.635 0.575 3.225 ;
        RECT 0.345 2.405 2.035 2.635 ;
        RECT 1.805 1.510 2.035 2.405 ;
        RECT 0.245 1.280 2.035 1.510 ;
        RECT 2.265 2.615 2.615 3.215 ;
        RECT 3.665 2.990 4.915 3.220 ;
        RECT 12.210 3.160 14.425 3.390 ;
        RECT 3.665 2.615 3.895 2.990 ;
        RECT 2.265 2.385 3.895 2.615 ;
        RECT 4.125 2.420 4.455 2.760 ;
        RECT 0.245 0.810 0.475 1.280 ;
        RECT 2.265 1.095 2.495 2.385 ;
        RECT 2.265 0.865 2.770 1.095 ;
        RECT 4.225 1.075 4.455 2.420 ;
        RECT 4.685 1.910 4.915 2.990 ;
        RECT 6.165 2.760 6.395 2.955 ;
        RECT 8.765 2.760 8.995 3.130 ;
        RECT 5.145 2.300 5.375 2.760 ;
        RECT 6.165 2.530 8.995 2.760 ;
        RECT 10.440 2.845 11.080 3.075 ;
        RECT 9.855 2.300 10.155 2.525 ;
        RECT 5.145 2.070 10.155 2.300 ;
        RECT 4.225 0.845 4.630 1.075 ;
        RECT 5.465 0.790 5.695 2.070 ;
        RECT 10.440 1.840 10.670 2.845 ;
        RECT 12.210 2.050 12.440 3.160 ;
        RECT 14.195 3.050 14.425 3.160 ;
        RECT 15.235 3.160 16.420 3.390 ;
        RECT 15.235 3.050 15.465 3.160 ;
        RECT 6.690 1.610 10.670 1.840 ;
        RECT 11.550 1.820 12.440 2.050 ;
        RECT 6.045 1.380 6.275 1.590 ;
        RECT 6.045 1.150 9.230 1.380 ;
        RECT 9.000 0.760 9.230 1.150 ;
        RECT 9.990 1.000 10.330 1.610 ;
        RECT 10.925 0.760 11.155 1.590 ;
        RECT 11.550 1.000 11.890 1.820 ;
        RECT 12.890 1.590 13.120 2.525 ;
        RECT 12.120 1.360 13.120 1.590 ;
        RECT 12.120 0.760 12.350 1.360 ;
        RECT 13.415 1.130 13.755 2.930 ;
        RECT 14.195 2.820 15.465 3.050 ;
        RECT 15.730 2.405 15.960 2.930 ;
        RECT 13.995 2.175 15.960 2.405 ;
        RECT 15.730 1.680 15.960 2.175 ;
        RECT 16.190 1.910 16.420 3.160 ;
        RECT 16.650 1.680 18.690 1.755 ;
        RECT 15.730 1.525 18.690 1.680 ;
        RECT 15.730 1.450 16.880 1.525 ;
        RECT 12.950 0.790 13.755 1.130 ;
        RECT 16.650 0.810 16.880 1.450 ;
        RECT 9.000 0.530 12.350 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
MACRO gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.400 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.606000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.890 1.770 3.920 2.150 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.429500 ;
    PORT
      LAYER Metal1 ;
        RECT 14.660 1.025 15.210 1.685 ;
        RECT 14.660 0.660 16.255 1.025 ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.675500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.280 1.770 1.570 2.150 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.111200 ;
    PORT
      LAYER Metal1 ;
        RECT 18.435 2.280 18.800 3.380 ;
        RECT 20.475 2.280 21.180 3.380 ;
        RECT 18.435 2.030 21.180 2.280 ;
        RECT 20.715 1.175 21.180 2.030 ;
        RECT 18.490 0.940 21.180 1.175 ;
        RECT 18.490 0.780 18.720 0.940 ;
        RECT 20.715 0.550 21.180 0.940 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 22.400 4.220 ;
        RECT 1.310 2.865 1.650 3.620 ;
        RECT 3.050 2.845 3.390 3.620 ;
        RECT 7.350 2.990 7.690 3.620 ;
        RECT 9.485 2.790 9.715 3.620 ;
        RECT 14.655 3.280 14.995 3.620 ;
        RECT 16.750 2.570 16.985 3.620 ;
        RECT 17.465 2.570 17.700 3.620 ;
        RECT 19.455 2.530 19.795 3.620 ;
        RECT 21.550 2.570 21.780 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.895 22.830 4.350 ;
        RECT -0.430 1.760 9.600 1.895 ;
        RECT 12.515 1.760 22.830 1.895 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 9.600 1.760 12.515 1.895 ;
        RECT -0.430 -0.430 22.830 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.655 1.050 ;
        RECT 3.170 0.300 3.510 1.075 ;
        RECT 8.430 0.300 8.770 0.915 ;
        RECT 14.070 0.300 14.300 1.130 ;
        RECT 17.315 0.300 17.655 0.640 ;
        RECT 19.555 0.300 19.895 0.710 ;
        RECT 21.850 0.300 22.080 0.765 ;
        RECT 0.000 -0.300 22.400 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 2.635 0.575 3.225 ;
        RECT 0.345 2.405 2.035 2.635 ;
        RECT 1.805 1.510 2.035 2.405 ;
        RECT 0.245 1.280 2.035 1.510 ;
        RECT 2.265 2.615 2.615 3.215 ;
        RECT 3.665 2.990 4.915 3.220 ;
        RECT 12.210 3.160 14.425 3.390 ;
        RECT 3.665 2.615 3.895 2.990 ;
        RECT 2.265 2.385 3.895 2.615 ;
        RECT 4.125 2.420 4.455 2.760 ;
        RECT 0.245 0.810 0.475 1.280 ;
        RECT 2.265 1.095 2.495 2.385 ;
        RECT 2.265 0.865 2.770 1.095 ;
        RECT 4.225 1.075 4.455 2.420 ;
        RECT 4.685 1.910 4.915 2.990 ;
        RECT 6.165 2.760 6.395 2.955 ;
        RECT 8.765 2.760 8.995 3.130 ;
        RECT 5.145 2.300 5.375 2.760 ;
        RECT 6.165 2.530 8.995 2.760 ;
        RECT 10.440 2.845 11.080 3.075 ;
        RECT 9.855 2.300 10.155 2.525 ;
        RECT 5.145 2.070 10.155 2.300 ;
        RECT 4.225 0.845 4.630 1.075 ;
        RECT 5.465 0.790 5.695 2.070 ;
        RECT 10.440 1.840 10.670 2.845 ;
        RECT 12.210 2.050 12.440 3.160 ;
        RECT 14.195 3.050 14.425 3.160 ;
        RECT 15.235 3.160 16.440 3.390 ;
        RECT 15.235 3.050 15.465 3.160 ;
        RECT 6.690 1.610 10.670 1.840 ;
        RECT 11.550 1.820 12.440 2.050 ;
        RECT 6.045 1.380 6.275 1.590 ;
        RECT 6.045 1.150 9.230 1.380 ;
        RECT 9.000 0.760 9.230 1.150 ;
        RECT 9.990 1.000 10.330 1.610 ;
        RECT 10.925 0.760 11.155 1.590 ;
        RECT 11.550 1.000 11.890 1.820 ;
        RECT 12.890 1.590 13.120 2.525 ;
        RECT 12.120 1.360 13.120 1.590 ;
        RECT 12.120 0.760 12.350 1.360 ;
        RECT 13.415 1.130 13.755 2.930 ;
        RECT 14.195 2.820 15.465 3.050 ;
        RECT 15.730 2.405 15.960 2.930 ;
        RECT 13.995 2.175 15.960 2.405 ;
        RECT 15.730 1.680 15.960 2.175 ;
        RECT 16.210 1.910 16.440 3.160 ;
        RECT 15.730 1.450 20.485 1.680 ;
        RECT 12.950 0.790 13.755 1.130 ;
        RECT 16.650 0.810 16.880 1.450 ;
        RECT 9.000 0.530 12.350 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
MACRO gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.840 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.401500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.890 1.770 3.960 2.150 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.209500 ;
    PORT
      LAYER Metal1 ;
        RECT 16.715 1.785 18.115 2.150 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.096000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.650 1.700 15.955 2.150 ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.675500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.280 1.770 1.575 2.130 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.893200 ;
    PORT
      LAYER Metal1 ;
        RECT 20.825 0.860 21.335 3.380 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 21.840 4.220 ;
        RECT 1.205 2.930 1.555 3.620 ;
        RECT 3.010 3.005 3.350 3.620 ;
        RECT 7.530 3.445 7.870 3.620 ;
        RECT 10.730 3.445 11.070 3.620 ;
        RECT 15.125 2.930 15.465 3.620 ;
        RECT 17.270 2.930 17.610 3.620 ;
        RECT 19.365 2.810 19.595 3.620 ;
        RECT 20.085 2.530 20.315 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.940 22.270 4.350 ;
        RECT -0.430 1.760 3.225 1.940 ;
        RECT 14.255 1.760 22.270 1.940 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 3.225 1.760 14.255 1.940 ;
        RECT -0.430 -0.430 22.270 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 1.050 ;
        RECT 3.510 0.300 3.850 1.150 ;
        RECT 8.850 0.300 9.190 0.915 ;
        RECT 17.170 0.300 17.510 1.075 ;
        RECT 19.925 0.300 20.155 0.765 ;
        RECT 0.000 -0.300 21.840 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.590 0.475 3.225 ;
        RECT 2.285 2.725 2.515 3.225 ;
        RECT 3.650 3.110 5.095 3.340 ;
        RECT 5.850 3.215 7.300 3.345 ;
        RECT 8.180 3.215 10.480 3.390 ;
        RECT 11.300 3.215 12.750 3.295 ;
        RECT 5.850 3.155 12.750 3.215 ;
        RECT 5.850 3.110 8.410 3.155 ;
        RECT 3.650 2.725 3.880 3.110 ;
        RECT 0.245 2.360 2.055 2.590 ;
        RECT 1.825 1.510 2.055 2.360 ;
        RECT 0.245 1.280 2.055 1.510 ;
        RECT 2.285 2.490 3.880 2.725 ;
        RECT 0.245 0.810 0.475 1.280 ;
        RECT 2.285 1.105 2.515 2.490 ;
        RECT 4.250 1.205 4.590 2.880 ;
        RECT 4.865 1.895 5.095 3.110 ;
        RECT 7.070 2.985 8.410 3.110 ;
        RECT 10.245 3.065 12.750 3.155 ;
        RECT 13.045 3.120 14.815 3.355 ;
        RECT 10.245 2.985 11.530 3.065 ;
        RECT 5.325 2.295 5.555 2.940 ;
        RECT 6.290 2.755 6.630 2.880 ;
        RECT 8.770 2.755 9.110 2.925 ;
        RECT 6.290 2.525 9.110 2.755 ;
        RECT 9.490 2.755 9.830 2.925 ;
        RECT 11.970 2.755 12.310 2.835 ;
        RECT 9.490 2.525 12.310 2.755 ;
        RECT 5.325 2.065 10.270 2.295 ;
        RECT 5.325 2.040 6.035 2.065 ;
        RECT 2.285 0.765 2.715 1.105 ;
        RECT 4.250 0.865 4.915 1.205 ;
        RECT 5.805 0.865 6.035 2.040 ;
        RECT 11.280 1.835 11.510 2.525 ;
        RECT 13.045 2.295 13.275 3.120 ;
        RECT 6.265 1.375 6.495 1.685 ;
        RECT 7.030 1.605 11.510 1.835 ;
        RECT 12.400 2.060 13.275 2.295 ;
        RECT 6.265 1.145 10.880 1.375 ;
        RECT 10.650 0.760 10.880 1.145 ;
        RECT 11.170 0.990 11.510 1.605 ;
        RECT 11.745 0.760 12.000 1.735 ;
        RECT 12.400 1.220 12.630 2.060 ;
        RECT 13.505 1.830 13.735 2.430 ;
        RECT 12.290 0.990 12.630 1.220 ;
        RECT 12.895 1.600 13.735 1.830 ;
        RECT 12.895 0.760 13.125 1.600 ;
        RECT 14.065 1.220 14.295 2.890 ;
        RECT 14.585 2.700 14.815 3.120 ;
        RECT 15.695 3.090 17.035 3.325 ;
        RECT 15.695 2.700 15.925 3.090 ;
        RECT 14.585 2.465 15.925 2.700 ;
        RECT 16.185 2.465 16.535 2.805 ;
        RECT 16.805 2.700 17.035 3.090 ;
        RECT 17.885 3.035 19.035 3.270 ;
        RECT 17.885 2.700 18.115 3.035 ;
        RECT 16.805 2.465 18.115 2.700 ;
        RECT 13.410 1.075 14.295 1.220 ;
        RECT 16.185 1.075 16.415 2.465 ;
        RECT 18.345 1.610 18.575 2.805 ;
        RECT 18.805 2.005 19.035 3.035 ;
        RECT 18.345 1.555 20.595 1.610 ;
        RECT 16.645 1.325 20.595 1.555 ;
        RECT 13.410 0.990 16.415 1.075 ;
        RECT 14.065 0.845 16.415 0.990 ;
        RECT 19.205 1.270 20.595 1.325 ;
        RECT 19.205 0.790 19.435 1.270 ;
        RECT 10.650 0.530 13.125 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1
MACRO gf180mcu_fd_sc_mcu7t5v0__dffrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffrsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.960 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.401500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.890 1.770 3.960 2.150 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.209500 ;
    PORT
      LAYER Metal1 ;
        RECT 16.715 1.785 18.115 2.150 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.096000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.650 1.700 15.955 2.150 ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.675500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.310 1.770 1.575 2.130 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.055600 ;
    PORT
      LAYER Metal1 ;
        RECT 21.100 2.330 21.755 3.380 ;
        RECT 21.370 1.090 21.755 2.330 ;
        RECT 20.990 0.860 21.755 1.090 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 22.960 4.220 ;
        RECT 1.205 2.930 1.555 3.620 ;
        RECT 3.010 3.005 3.350 3.620 ;
        RECT 7.530 3.445 7.870 3.620 ;
        RECT 10.730 3.445 11.070 3.620 ;
        RECT 15.125 2.930 15.465 3.620 ;
        RECT 17.270 2.930 17.610 3.620 ;
        RECT 19.365 2.810 19.595 3.620 ;
        RECT 20.085 2.570 20.315 3.620 ;
        RECT 22.125 2.570 22.355 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.940 23.390 4.350 ;
        RECT -0.430 1.760 3.225 1.940 ;
        RECT 14.255 1.760 23.390 1.940 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 3.225 1.760 14.255 1.940 ;
        RECT -0.430 -0.430 23.390 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 1.050 ;
        RECT 3.510 0.300 3.850 1.150 ;
        RECT 8.850 0.300 9.190 0.915 ;
        RECT 17.170 0.300 17.510 1.075 ;
        RECT 19.925 0.300 20.155 0.765 ;
        RECT 22.210 0.300 22.550 0.640 ;
        RECT 0.000 -0.300 22.960 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.590 0.475 3.225 ;
        RECT 2.285 2.725 2.515 3.225 ;
        RECT 3.650 3.110 5.095 3.340 ;
        RECT 5.850 3.215 7.300 3.345 ;
        RECT 8.180 3.215 10.480 3.390 ;
        RECT 11.300 3.215 12.750 3.295 ;
        RECT 5.850 3.155 12.750 3.215 ;
        RECT 5.850 3.110 8.410 3.155 ;
        RECT 3.650 2.725 3.880 3.110 ;
        RECT 0.245 2.360 2.055 2.590 ;
        RECT 1.825 1.510 2.055 2.360 ;
        RECT 0.245 1.280 2.055 1.510 ;
        RECT 2.285 2.490 3.880 2.725 ;
        RECT 0.245 0.810 0.475 1.280 ;
        RECT 2.285 1.105 2.515 2.490 ;
        RECT 4.250 1.205 4.590 2.880 ;
        RECT 4.865 1.895 5.095 3.110 ;
        RECT 7.070 2.985 8.410 3.110 ;
        RECT 10.245 3.065 12.750 3.155 ;
        RECT 13.045 3.120 14.815 3.355 ;
        RECT 10.245 2.985 11.530 3.065 ;
        RECT 5.325 2.295 5.555 2.940 ;
        RECT 6.290 2.755 6.630 2.880 ;
        RECT 8.770 2.755 9.110 2.925 ;
        RECT 6.290 2.525 9.110 2.755 ;
        RECT 9.490 2.755 9.830 2.925 ;
        RECT 11.970 2.755 12.310 2.835 ;
        RECT 9.490 2.525 12.310 2.755 ;
        RECT 5.325 2.065 10.270 2.295 ;
        RECT 5.325 2.040 6.035 2.065 ;
        RECT 2.285 0.765 2.715 1.105 ;
        RECT 4.250 0.865 4.915 1.205 ;
        RECT 5.805 0.865 6.035 2.040 ;
        RECT 11.280 1.835 11.510 2.525 ;
        RECT 13.045 2.295 13.275 3.120 ;
        RECT 6.265 1.375 6.495 1.685 ;
        RECT 7.030 1.605 11.510 1.835 ;
        RECT 12.400 2.060 13.275 2.295 ;
        RECT 6.265 1.145 10.880 1.375 ;
        RECT 10.650 0.760 10.880 1.145 ;
        RECT 11.170 0.990 11.510 1.605 ;
        RECT 11.745 0.760 12.000 1.735 ;
        RECT 12.400 1.220 12.630 2.060 ;
        RECT 13.505 1.830 13.735 2.430 ;
        RECT 12.290 0.990 12.630 1.220 ;
        RECT 12.895 1.600 13.735 1.830 ;
        RECT 12.895 0.760 13.125 1.600 ;
        RECT 14.065 1.220 14.295 2.890 ;
        RECT 14.585 2.700 14.815 3.120 ;
        RECT 15.695 3.090 17.035 3.325 ;
        RECT 15.695 2.700 15.925 3.090 ;
        RECT 14.585 2.465 15.925 2.700 ;
        RECT 16.185 2.465 16.535 2.805 ;
        RECT 16.805 2.700 17.035 3.090 ;
        RECT 17.885 3.035 19.035 3.270 ;
        RECT 17.885 2.700 18.115 3.035 ;
        RECT 16.805 2.465 18.115 2.700 ;
        RECT 13.410 1.075 14.295 1.220 ;
        RECT 16.185 1.075 16.415 2.465 ;
        RECT 18.345 1.555 18.575 2.805 ;
        RECT 18.805 2.005 19.035 3.035 ;
        RECT 20.305 1.555 21.120 1.755 ;
        RECT 16.645 1.525 21.120 1.555 ;
        RECT 16.645 1.325 20.595 1.525 ;
        RECT 13.410 0.990 16.415 1.075 ;
        RECT 14.065 0.845 16.415 0.990 ;
        RECT 19.205 0.790 19.435 1.325 ;
        RECT 10.650 0.530 13.125 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffrsnq_2
MACRO gf180mcu_fd_sc_mcu7t5v0__dffrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffrsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.200 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.456500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.850 1.650 3.960 2.150 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.177000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.715 1.785 18.115 2.130 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.096000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.565 1.670 15.955 2.225 ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.675500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 0.600 1.070 2.150 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.111200 ;
    PORT
      LAYER Metal1 ;
        RECT 21.045 2.360 21.335 3.380 ;
        RECT 23.060 2.360 23.420 3.380 ;
        RECT 21.045 2.280 23.420 2.360 ;
        RECT 21.045 2.125 24.005 2.280 ;
        RECT 23.140 1.315 24.005 2.125 ;
        RECT 21.045 1.085 24.005 1.315 ;
        RECT 21.045 0.655 21.275 1.085 ;
        RECT 23.140 0.600 24.005 1.085 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 25.200 4.220 ;
        RECT 1.205 2.930 1.555 3.620 ;
        RECT 3.010 3.005 3.350 3.620 ;
        RECT 7.530 3.445 7.870 3.620 ;
        RECT 10.730 3.445 11.070 3.620 ;
        RECT 15.125 2.930 15.465 3.620 ;
        RECT 17.270 2.930 17.610 3.620 ;
        RECT 19.365 2.730 19.595 3.620 ;
        RECT 20.085 2.530 20.315 3.620 ;
        RECT 22.070 2.620 22.410 3.620 ;
        RECT 24.165 2.530 24.395 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 25.630 4.350 ;
        RECT -0.430 1.760 3.225 1.885 ;
        RECT 14.255 1.760 25.630 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 3.225 1.760 14.255 1.885 ;
        RECT -0.430 -0.430 25.630 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 1.160 ;
        RECT 3.510 0.300 3.850 1.150 ;
        RECT 8.850 0.300 9.190 0.915 ;
        RECT 17.170 0.300 17.510 1.075 ;
        RECT 19.925 0.300 20.155 0.905 ;
        RECT 22.165 0.300 22.395 0.765 ;
        RECT 24.405 0.300 24.635 0.905 ;
        RECT 0.000 -0.300 25.200 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.700 0.475 3.225 ;
        RECT 2.285 2.725 2.515 3.225 ;
        RECT 3.650 3.160 4.995 3.390 ;
        RECT 5.780 3.215 7.300 3.390 ;
        RECT 8.180 3.215 10.480 3.390 ;
        RECT 11.300 3.215 12.750 3.295 ;
        RECT 5.780 3.160 12.750 3.215 ;
        RECT 3.650 2.725 3.880 3.160 ;
        RECT 0.245 2.380 2.035 2.700 ;
        RECT 0.245 0.810 0.475 2.380 ;
        RECT 1.805 1.280 2.035 2.380 ;
        RECT 2.285 2.490 3.880 2.725 ;
        RECT 2.285 1.105 2.515 2.490 ;
        RECT 4.305 1.205 4.535 2.930 ;
        RECT 4.765 1.895 4.995 3.160 ;
        RECT 7.070 2.985 8.410 3.160 ;
        RECT 10.245 3.065 12.750 3.160 ;
        RECT 13.045 3.120 14.815 3.355 ;
        RECT 10.245 2.985 11.530 3.065 ;
        RECT 5.325 2.295 5.555 2.940 ;
        RECT 6.290 2.755 6.630 2.885 ;
        RECT 8.770 2.755 9.110 2.930 ;
        RECT 6.290 2.525 9.110 2.755 ;
        RECT 9.490 2.755 9.830 2.930 ;
        RECT 11.970 2.755 12.310 2.835 ;
        RECT 9.490 2.525 12.310 2.755 ;
        RECT 5.325 2.065 10.360 2.295 ;
        RECT 5.325 2.040 6.035 2.065 ;
        RECT 2.285 0.765 2.715 1.105 ;
        RECT 4.305 0.865 4.915 1.205 ;
        RECT 5.805 0.865 6.035 2.040 ;
        RECT 11.280 1.835 11.510 2.525 ;
        RECT 13.045 2.295 13.275 3.120 ;
        RECT 6.265 1.375 6.495 1.685 ;
        RECT 7.030 1.605 11.510 1.835 ;
        RECT 12.400 2.060 13.275 2.295 ;
        RECT 6.265 1.145 10.880 1.375 ;
        RECT 10.650 0.760 10.880 1.145 ;
        RECT 11.170 0.990 11.510 1.605 ;
        RECT 11.745 0.760 12.000 1.735 ;
        RECT 12.400 1.220 12.630 2.060 ;
        RECT 13.505 1.830 13.735 2.430 ;
        RECT 12.290 0.990 12.630 1.220 ;
        RECT 12.895 1.600 13.735 1.830 ;
        RECT 12.895 0.760 13.125 1.600 ;
        RECT 14.065 1.220 14.295 2.890 ;
        RECT 14.585 2.700 14.815 3.120 ;
        RECT 15.695 3.090 17.035 3.325 ;
        RECT 15.695 2.700 15.925 3.090 ;
        RECT 14.585 2.465 15.925 2.700 ;
        RECT 16.185 2.465 16.535 2.805 ;
        RECT 16.805 2.700 17.035 3.090 ;
        RECT 17.885 3.035 19.035 3.270 ;
        RECT 17.885 2.700 18.115 3.035 ;
        RECT 16.805 2.465 18.115 2.700 ;
        RECT 13.410 1.075 14.295 1.220 ;
        RECT 16.185 1.075 16.415 2.465 ;
        RECT 18.345 1.555 18.575 2.805 ;
        RECT 18.805 2.005 19.035 3.035 ;
        RECT 20.305 1.555 22.890 1.785 ;
        RECT 16.645 1.325 20.595 1.555 ;
        RECT 13.410 0.990 16.415 1.075 ;
        RECT 14.065 0.845 16.415 0.990 ;
        RECT 19.205 0.790 19.435 1.325 ;
        RECT 10.650 0.530 13.125 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffrsnq_4
MACRO gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.160 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.468500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.890 1.770 4.030 2.150 ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.141500 ;
    PORT
      LAYER Metal1 ;
        RECT 14.090 1.770 15.285 2.150 ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.675500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.280 1.765 1.590 2.130 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.014700 ;
    PORT
      LAYER Metal1 ;
        RECT 19.045 2.190 19.815 3.380 ;
        RECT 19.425 1.160 19.815 2.190 ;
        RECT 19.300 0.550 19.815 1.160 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 20.160 4.220 ;
        RECT 1.310 2.930 1.650 3.620 ;
        RECT 3.240 2.845 3.580 3.620 ;
        RECT 7.675 3.445 8.015 3.620 ;
        RECT 10.275 3.005 10.615 3.620 ;
        RECT 14.295 3.005 14.635 3.620 ;
        RECT 16.710 2.530 16.940 3.620 ;
        RECT 18.450 2.530 18.680 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 20.590 4.350 ;
        RECT -0.430 1.760 9.135 1.885 ;
        RECT 15.165 1.760 20.590 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 9.135 1.760 15.165 1.885 ;
        RECT -0.430 -0.430 20.590 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 1.050 ;
        RECT 3.150 0.300 3.490 1.075 ;
        RECT 7.455 0.300 7.795 1.075 ;
        RECT 16.555 0.300 16.895 1.050 ;
        RECT 18.450 0.300 18.680 0.765 ;
        RECT 0.000 -0.300 20.160 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 2.595 0.575 3.225 ;
        RECT 2.385 2.615 2.615 3.225 ;
        RECT 3.810 3.160 5.115 3.390 ;
        RECT 8.270 3.215 9.915 3.390 ;
        RECT 3.810 2.615 4.040 3.160 ;
        RECT 0.345 2.360 2.090 2.595 ;
        RECT 1.860 1.510 2.090 2.360 ;
        RECT 0.245 1.280 2.090 1.510 ;
        RECT 2.385 2.380 4.040 2.615 ;
        RECT 0.245 0.810 0.475 1.280 ;
        RECT 2.385 1.150 2.620 2.380 ;
        RECT 2.385 0.810 2.715 1.150 ;
        RECT 4.270 0.790 4.610 2.930 ;
        RECT 4.885 1.930 5.115 3.160 ;
        RECT 6.115 3.160 9.915 3.215 ;
        RECT 6.115 2.985 8.500 3.160 ;
        RECT 5.345 1.995 5.575 2.985 ;
        RECT 6.115 2.240 6.455 2.985 ;
        RECT 9.035 2.455 9.375 2.930 ;
        RECT 9.685 2.775 9.915 3.160 ;
        RECT 10.845 3.065 12.315 3.295 ;
        RECT 10.845 2.775 11.075 3.065 ;
        RECT 9.685 2.540 11.075 2.775 ;
        RECT 7.015 2.310 9.375 2.455 ;
        RECT 11.305 2.310 11.645 2.780 ;
        RECT 7.015 2.225 11.645 2.310 ;
        RECT 9.035 2.080 11.645 2.225 ;
        RECT 11.930 2.550 12.895 2.780 ;
        RECT 13.630 2.775 13.860 2.845 ;
        RECT 15.370 2.775 15.600 2.885 ;
        RECT 5.345 1.765 8.235 1.995 ;
        RECT 5.345 0.790 5.675 1.765 ;
        RECT 6.000 1.305 8.340 1.535 ;
        RECT 8.110 0.760 8.340 1.305 ;
        RECT 9.875 0.990 10.215 2.080 ;
        RECT 10.810 0.760 11.040 1.615 ;
        RECT 11.930 1.130 12.160 2.550 ;
        RECT 13.630 2.540 15.600 2.775 ;
        RECT 13.630 1.220 13.860 2.540 ;
        RECT 17.730 2.105 17.960 3.380 ;
        RECT 15.755 1.860 17.960 2.105 ;
        RECT 17.730 1.840 17.960 1.860 ;
        RECT 15.880 1.395 17.335 1.630 ;
        RECT 17.730 1.500 19.120 1.840 ;
        RECT 11.270 0.790 12.160 1.130 ;
        RECT 12.555 0.990 14.495 1.220 ;
        RECT 8.110 0.530 11.040 0.760 ;
        RECT 11.930 0.760 12.160 0.790 ;
        RECT 15.880 0.760 16.110 1.395 ;
        RECT 17.730 0.805 17.960 1.500 ;
        RECT 11.930 0.530 16.110 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
MACRO gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.468500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.890 1.770 4.030 2.150 ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.141500 ;
    PORT
      LAYER Metal1 ;
        RECT 14.090 1.770 15.285 2.150 ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.675500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 1.765 1.590 2.130 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.298600 ;
    PORT
      LAYER Metal1 ;
        RECT 19.530 2.330 20.370 3.380 ;
        RECT 19.950 1.020 20.370 2.330 ;
        RECT 19.330 0.550 20.370 1.020 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 21.280 4.220 ;
        RECT 1.310 2.930 1.650 3.620 ;
        RECT 3.240 2.845 3.580 3.620 ;
        RECT 7.675 3.445 8.015 3.620 ;
        RECT 10.275 3.005 10.615 3.620 ;
        RECT 14.295 3.005 14.635 3.620 ;
        RECT 16.810 2.530 17.040 3.620 ;
        RECT 18.550 2.530 18.780 3.620 ;
        RECT 20.790 2.530 21.020 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 21.710 4.350 ;
        RECT -0.430 1.760 9.135 1.885 ;
        RECT 15.165 1.760 21.710 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 9.135 1.760 15.165 1.885 ;
        RECT -0.430 -0.430 21.710 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 1.050 ;
        RECT 3.150 0.300 3.490 1.075 ;
        RECT 7.455 0.300 7.795 1.075 ;
        RECT 16.555 0.300 16.895 0.835 ;
        RECT 18.550 0.300 18.780 0.890 ;
        RECT 20.790 0.300 21.020 0.890 ;
        RECT 0.000 -0.300 21.280 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 2.595 0.575 3.225 ;
        RECT 2.385 2.615 2.615 3.225 ;
        RECT 3.810 3.160 5.115 3.390 ;
        RECT 8.270 3.215 9.915 3.390 ;
        RECT 3.810 2.615 4.040 3.160 ;
        RECT 0.345 2.360 2.090 2.595 ;
        RECT 1.860 1.510 2.090 2.360 ;
        RECT 0.245 1.280 2.090 1.510 ;
        RECT 2.385 2.380 4.040 2.615 ;
        RECT 0.245 0.810 0.475 1.280 ;
        RECT 2.385 1.150 2.620 2.380 ;
        RECT 2.385 0.810 2.715 1.150 ;
        RECT 4.270 0.790 4.610 2.930 ;
        RECT 4.885 1.930 5.115 3.160 ;
        RECT 6.115 3.160 9.915 3.215 ;
        RECT 6.115 2.985 8.500 3.160 ;
        RECT 5.345 1.995 5.575 2.985 ;
        RECT 6.115 2.240 6.455 2.985 ;
        RECT 9.035 2.455 9.375 2.930 ;
        RECT 9.685 2.775 9.915 3.160 ;
        RECT 10.845 3.065 12.315 3.295 ;
        RECT 10.845 2.775 11.075 3.065 ;
        RECT 9.685 2.540 11.075 2.775 ;
        RECT 7.015 2.310 9.375 2.455 ;
        RECT 11.305 2.310 11.645 2.780 ;
        RECT 7.015 2.225 11.645 2.310 ;
        RECT 9.035 2.080 11.645 2.225 ;
        RECT 11.930 2.550 12.895 2.780 ;
        RECT 13.630 2.775 13.860 2.845 ;
        RECT 15.370 2.775 15.600 2.885 ;
        RECT 5.345 1.765 8.235 1.995 ;
        RECT 5.345 0.790 5.675 1.765 ;
        RECT 6.000 1.305 8.340 1.535 ;
        RECT 8.110 0.760 8.340 1.305 ;
        RECT 9.875 0.990 10.215 2.080 ;
        RECT 10.810 0.760 11.040 1.615 ;
        RECT 11.930 1.130 12.160 2.550 ;
        RECT 13.630 2.540 15.600 2.775 ;
        RECT 13.630 1.220 13.860 2.540 ;
        RECT 17.830 2.105 18.060 3.380 ;
        RECT 15.755 1.860 18.060 2.105 ;
        RECT 17.730 1.840 18.060 1.860 ;
        RECT 15.880 1.395 17.335 1.630 ;
        RECT 17.730 1.500 19.690 1.840 ;
        RECT 11.270 0.790 12.160 1.130 ;
        RECT 12.555 0.990 14.495 1.220 ;
        RECT 8.110 0.530 11.040 0.760 ;
        RECT 11.930 0.760 12.160 0.790 ;
        RECT 15.880 0.760 16.110 1.395 ;
        RECT 11.930 0.530 16.110 0.760 ;
        RECT 17.730 0.550 17.960 1.500 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
MACRO gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.080 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.468500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.890 1.770 4.030 2.150 ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.141500 ;
    PORT
      LAYER Metal1 ;
        RECT 14.090 1.770 15.285 2.150 ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.675500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.280 1.765 1.590 2.130 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.597200 ;
    PORT
      LAYER Metal1 ;
        RECT 20.050 2.290 20.280 3.380 ;
        RECT 21.670 2.290 22.535 3.380 ;
        RECT 20.050 2.060 22.535 2.290 ;
        RECT 22.010 1.315 22.535 2.060 ;
        RECT 20.045 1.085 22.535 1.315 ;
        RECT 20.045 0.550 20.280 1.085 ;
        RECT 22.010 0.550 22.535 1.085 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 24.080 4.220 ;
        RECT 1.310 2.930 1.650 3.620 ;
        RECT 3.240 2.845 3.580 3.620 ;
        RECT 7.675 3.445 8.015 3.620 ;
        RECT 10.275 3.005 10.615 3.620 ;
        RECT 14.295 3.005 14.635 3.620 ;
        RECT 16.705 2.530 16.935 3.620 ;
        RECT 18.750 2.530 18.980 3.620 ;
        RECT 21.170 2.530 21.400 3.620 ;
        RECT 23.410 2.530 23.640 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 24.510 4.350 ;
        RECT -0.430 1.760 9.135 1.885 ;
        RECT 15.165 1.760 24.510 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 9.135 1.760 15.165 1.885 ;
        RECT -0.430 -0.430 24.510 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 1.050 ;
        RECT 3.150 0.300 3.490 1.075 ;
        RECT 7.455 0.300 7.795 1.075 ;
        RECT 16.555 0.300 16.895 0.835 ;
        RECT 18.850 0.300 19.080 0.890 ;
        RECT 21.115 0.300 21.455 0.835 ;
        RECT 23.410 0.300 23.640 0.890 ;
        RECT 0.000 -0.300 24.080 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 2.595 0.575 3.225 ;
        RECT 2.385 2.615 2.615 3.225 ;
        RECT 3.810 3.160 5.115 3.390 ;
        RECT 8.270 3.215 9.915 3.390 ;
        RECT 3.810 2.615 4.040 3.160 ;
        RECT 0.345 2.360 2.090 2.595 ;
        RECT 1.860 1.510 2.090 2.360 ;
        RECT 0.245 1.280 2.090 1.510 ;
        RECT 2.385 2.380 4.040 2.615 ;
        RECT 0.245 0.810 0.475 1.280 ;
        RECT 2.385 1.150 2.620 2.380 ;
        RECT 2.385 0.810 2.715 1.150 ;
        RECT 4.270 0.790 4.610 2.930 ;
        RECT 4.885 1.930 5.115 3.160 ;
        RECT 6.115 3.160 9.915 3.215 ;
        RECT 6.115 2.985 8.500 3.160 ;
        RECT 5.345 1.995 5.575 2.985 ;
        RECT 6.115 2.240 6.455 2.985 ;
        RECT 9.035 2.455 9.375 2.930 ;
        RECT 9.685 2.775 9.915 3.160 ;
        RECT 10.845 3.065 12.315 3.295 ;
        RECT 10.845 2.775 11.075 3.065 ;
        RECT 9.685 2.540 11.075 2.775 ;
        RECT 7.015 2.310 9.375 2.455 ;
        RECT 11.305 2.310 11.645 2.780 ;
        RECT 7.015 2.225 11.645 2.310 ;
        RECT 9.035 2.080 11.645 2.225 ;
        RECT 11.930 2.550 12.895 2.780 ;
        RECT 13.630 2.775 13.860 2.845 ;
        RECT 15.370 2.775 15.600 2.885 ;
        RECT 5.345 1.765 8.235 1.995 ;
        RECT 5.345 0.790 5.675 1.765 ;
        RECT 6.000 1.305 8.340 1.535 ;
        RECT 8.110 0.760 8.340 1.305 ;
        RECT 9.875 0.990 10.215 2.080 ;
        RECT 10.810 0.760 11.040 1.615 ;
        RECT 11.930 1.130 12.160 2.550 ;
        RECT 13.630 2.540 15.600 2.775 ;
        RECT 13.630 1.220 13.860 2.540 ;
        RECT 17.730 2.105 17.960 3.380 ;
        RECT 15.755 1.860 17.960 2.105 ;
        RECT 17.730 1.785 17.960 1.860 ;
        RECT 15.880 1.395 17.335 1.630 ;
        RECT 17.730 1.555 21.605 1.785 ;
        RECT 11.270 0.790 12.160 1.130 ;
        RECT 12.555 0.990 14.495 1.220 ;
        RECT 8.110 0.530 11.040 0.760 ;
        RECT 11.930 0.760 12.160 0.790 ;
        RECT 15.880 0.760 16.110 1.395 ;
        RECT 11.930 0.530 16.110 0.760 ;
        RECT 17.730 0.550 17.960 1.555 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
MACRO gf180mcu_fd_sc_mcu7t5v0__dlya_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlya_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.160 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 1.210 1.845 1.610 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 5.650 0.550 6.020 3.380 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 6.160 4.220 ;
        RECT 1.210 2.540 1.550 3.620 ;
        RECT 4.645 2.530 4.875 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 6.590 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.590 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 0.980 ;
        RECT 4.545 0.300 4.775 0.690 ;
        RECT 0.000 -0.300 6.160 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.255 0.475 2.825 ;
        RECT 0.245 2.025 2.135 2.255 ;
        RECT 0.245 0.640 0.475 2.025 ;
        RECT 2.385 1.725 2.615 2.825 ;
        RECT 3.105 2.280 3.335 2.710 ;
        RECT 3.105 2.050 5.215 2.280 ;
        RECT 2.385 1.495 4.180 1.725 ;
        RECT 2.385 0.640 2.715 1.495 ;
        RECT 4.985 1.180 5.215 2.050 ;
        RECT 3.870 0.950 5.215 1.180 ;
        RECT 3.870 0.765 4.105 0.950 ;
        RECT 3.145 0.530 4.105 0.765 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlya_1
MACRO gf180mcu_fd_sc_mcu7t5v0__dlya_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlya_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 1.210 1.590 1.610 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.188900 ;
    PORT
      LAYER Metal1 ;
        RECT 5.660 0.805 6.070 3.380 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.280 4.220 ;
        RECT 1.210 2.540 1.550 3.620 ;
        RECT 4.640 2.530 4.870 3.620 ;
        RECT 6.785 2.530 7.020 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 7.710 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 0.980 ;
        RECT 4.545 0.300 4.775 0.690 ;
        RECT 6.785 0.300 7.015 1.145 ;
        RECT 0.000 -0.300 7.280 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.310 0.475 2.825 ;
        RECT 0.245 2.075 2.035 2.310 ;
        RECT 0.245 0.640 0.475 2.075 ;
        RECT 1.805 1.970 2.035 2.075 ;
        RECT 2.385 1.790 2.615 2.825 ;
        RECT 3.105 2.280 3.335 2.710 ;
        RECT 3.105 2.050 5.375 2.280 ;
        RECT 2.385 1.550 4.055 1.790 ;
        RECT 2.385 0.640 2.715 1.550 ;
        RECT 5.145 1.250 5.375 2.050 ;
        RECT 4.050 1.020 5.375 1.250 ;
        RECT 4.050 0.765 4.285 1.020 ;
        RECT 3.145 0.530 4.285 0.765 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlya_2
MACRO gf180mcu_fd_sc_mcu7t5v0__dlya_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlya_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.210 2.150 1.590 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal1 ;
        RECT 5.680 2.580 5.910 3.160 ;
        RECT 7.820 2.580 8.390 3.160 ;
        RECT 5.680 2.350 8.390 2.580 ;
        RECT 7.820 1.405 8.390 2.350 ;
        RECT 5.630 1.170 8.390 1.405 ;
        RECT 5.630 0.600 5.860 1.170 ;
        RECT 7.870 0.600 8.390 1.170 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 9.520 4.220 ;
        RECT 1.270 2.635 1.500 3.620 ;
        RECT 4.455 2.660 4.795 3.620 ;
        RECT 6.645 2.810 6.985 3.620 ;
        RECT 8.890 2.605 9.120 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 9.950 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.315 0.300 1.655 0.845 ;
        RECT 4.330 0.300 4.560 0.905 ;
        RECT 6.750 0.300 6.980 0.940 ;
        RECT 8.990 0.300 9.220 0.940 ;
        RECT 0.000 -0.300 9.520 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.250 2.405 0.480 2.980 ;
        RECT 2.390 2.640 2.720 2.980 ;
        RECT 0.250 2.175 2.095 2.405 ;
        RECT 0.250 0.560 0.480 2.175 ;
        RECT 2.490 1.830 2.720 2.640 ;
        RECT 3.260 2.295 3.490 2.980 ;
        RECT 3.260 2.060 4.445 2.295 ;
        RECT 4.215 2.025 4.445 2.060 ;
        RECT 2.490 1.600 3.985 1.830 ;
        RECT 4.215 1.685 7.060 2.025 ;
        RECT 2.490 0.560 2.720 1.600 ;
        RECT 4.215 1.370 4.445 1.685 ;
        RECT 3.210 1.135 4.445 1.370 ;
        RECT 3.210 0.560 3.440 1.135 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlya_4
MACRO gf180mcu_fd_sc_mcu7t5v0__dlyb_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlyb_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.960 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.930 1.200 3.355 1.600 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 8.215 2.710 8.600 3.195 ;
        RECT 6.810 2.330 8.600 2.710 ;
        RECT 8.370 0.675 8.600 2.330 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 8.960 4.220 ;
        RECT 1.485 3.285 1.825 3.620 ;
        RECT 6.565 3.175 6.905 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 9.390 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.390 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.585 0.300 1.925 0.635 ;
        RECT 6.720 0.300 6.950 0.690 ;
        RECT 0.000 -0.300 8.960 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.405 0.585 3.105 ;
        RECT 0.245 2.065 3.265 2.405 ;
        RECT 0.245 0.900 0.475 2.065 ;
        RECT 3.720 1.910 3.950 3.160 ;
        RECT 4.540 2.465 4.770 3.160 ;
        RECT 4.540 2.235 6.155 2.465 ;
        RECT 3.720 1.680 5.485 1.910 ;
        RECT 0.245 0.670 0.585 0.900 ;
        RECT 3.720 0.770 4.105 1.680 ;
        RECT 5.835 1.625 6.155 2.235 ;
        RECT 5.835 1.395 7.975 1.625 ;
        RECT 5.835 1.055 6.155 1.395 ;
        RECT 4.540 0.715 6.155 1.055 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlyb_1
MACRO gf180mcu_fd_sc_mcu7t5v0__dlyb_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlyb_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.930 1.200 3.355 1.600 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.060800 ;
    PORT
      LAYER Metal1 ;
        RECT 8.420 2.340 8.860 3.390 ;
        RECT 8.420 2.105 9.380 2.340 ;
        RECT 8.930 1.215 9.380 2.105 ;
        RECT 8.370 0.960 9.380 1.215 ;
        RECT 8.370 0.530 8.600 0.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 10.080 4.220 ;
        RECT 1.485 3.285 1.825 3.620 ;
        RECT 6.565 3.175 7.685 3.620 ;
        RECT 7.345 2.530 7.685 3.175 ;
        RECT 9.435 2.570 9.775 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 10.510 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.585 0.300 1.925 0.635 ;
        RECT 6.720 0.300 6.950 0.690 ;
        RECT 9.435 0.300 9.775 0.635 ;
        RECT 0.000 -0.300 10.080 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.405 0.585 3.105 ;
        RECT 0.245 2.065 3.265 2.405 ;
        RECT 0.245 0.900 0.475 2.065 ;
        RECT 3.720 1.910 3.950 3.160 ;
        RECT 4.540 2.465 4.770 3.160 ;
        RECT 4.540 2.235 6.155 2.465 ;
        RECT 3.720 1.680 5.485 1.910 ;
        RECT 5.835 1.855 6.155 2.235 ;
        RECT 0.245 0.670 0.585 0.900 ;
        RECT 3.720 0.770 4.105 1.680 ;
        RECT 5.835 1.625 8.540 1.855 ;
        RECT 5.835 1.055 6.155 1.625 ;
        RECT 4.540 0.715 6.155 1.055 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlyb_2
MACRO gf180mcu_fd_sc_mcu7t5v0__dlyb_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlyb_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.320 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.930 1.200 3.360 1.600 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.304600 ;
    PORT
      LAYER Metal1 ;
        RECT 8.420 2.340 8.650 3.380 ;
        RECT 10.610 2.340 11.180 3.380 ;
        RECT 8.420 2.105 11.180 2.340 ;
        RECT 10.610 1.215 11.180 2.105 ;
        RECT 8.370 0.960 11.180 1.215 ;
        RECT 8.370 0.530 8.600 0.960 ;
        RECT 10.610 0.550 11.180 0.960 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 12.320 4.220 ;
        RECT 1.485 3.285 1.825 3.620 ;
        RECT 6.565 3.175 7.685 3.620 ;
        RECT 7.355 2.530 7.685 3.175 ;
        RECT 9.440 2.570 9.670 3.620 ;
        RECT 11.630 2.530 11.860 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 12.750 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.750 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.585 0.300 1.925 0.635 ;
        RECT 6.720 0.300 6.950 0.690 ;
        RECT 9.435 0.300 9.775 0.635 ;
        RECT 11.730 0.300 11.960 1.115 ;
        RECT 0.000 -0.300 12.320 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.405 0.585 3.105 ;
        RECT 0.245 2.065 3.265 2.405 ;
        RECT 0.245 0.900 0.475 2.065 ;
        RECT 3.720 1.910 3.950 3.160 ;
        RECT 4.540 2.465 4.770 3.160 ;
        RECT 4.540 2.235 6.155 2.465 ;
        RECT 3.720 1.680 5.485 1.910 ;
        RECT 5.835 1.855 6.155 2.235 ;
        RECT 0.245 0.670 0.585 0.900 ;
        RECT 3.720 0.770 4.105 1.680 ;
        RECT 5.835 1.625 10.360 1.855 ;
        RECT 5.835 1.055 6.155 1.625 ;
        RECT 4.540 0.715 6.155 1.055 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlyb_4
MACRO gf180mcu_fd_sc_mcu7t5v0__dlyc_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlyc_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.000 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.905 1.200 3.330 1.600 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 13.370 2.710 13.755 3.195 ;
        RECT 11.965 2.330 13.755 2.710 ;
        RECT 13.525 0.675 13.755 2.330 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 14.000 4.220 ;
        RECT 1.460 3.285 1.800 3.620 ;
        RECT 6.440 3.285 6.780 3.620 ;
        RECT 11.720 3.175 12.060 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 14.430 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.430 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.560 0.300 1.900 0.635 ;
        RECT 6.640 0.300 6.980 0.635 ;
        RECT 12.115 0.300 12.345 0.690 ;
        RECT 0.000 -0.300 14.000 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.220 2.405 0.560 3.105 ;
        RECT 0.220 2.065 3.240 2.405 ;
        RECT 0.220 0.670 0.560 2.065 ;
        RECT 3.695 1.805 3.925 3.160 ;
        RECT 4.360 2.875 5.765 3.105 ;
        RECT 3.695 1.465 5.305 1.805 ;
        RECT 5.535 1.750 5.765 2.875 ;
        RECT 8.875 1.965 9.260 3.160 ;
        RECT 9.695 2.465 9.925 3.160 ;
        RECT 9.695 2.235 11.665 2.465 ;
        RECT 5.535 1.520 8.090 1.750 ;
        RECT 8.875 1.535 11.055 1.965 ;
        RECT 11.345 1.625 11.665 2.235 ;
        RECT 3.695 0.770 4.080 1.465 ;
        RECT 5.535 1.000 5.765 1.520 ;
        RECT 4.460 0.770 5.765 1.000 ;
        RECT 8.875 0.715 9.105 1.535 ;
        RECT 11.345 1.395 13.130 1.625 ;
        RECT 11.345 1.055 11.665 1.395 ;
        RECT 9.695 0.715 11.665 1.055 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlyc_1
MACRO gf180mcu_fd_sc_mcu7t5v0__dlyc_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlyc_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.120 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.930 1.200 3.350 1.600 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.281700 ;
    PORT
      LAYER Metal1 ;
        RECT 13.395 0.675 13.910 3.195 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 15.120 4.220 ;
        RECT 1.485 3.285 1.825 3.620 ;
        RECT 6.465 3.285 6.805 3.620 ;
        RECT 11.745 3.175 12.085 3.620 ;
        RECT 14.465 2.705 14.805 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 15.550 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 15.550 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.585 0.300 1.925 0.635 ;
        RECT 6.665 0.300 7.005 0.635 ;
        RECT 11.925 0.300 12.155 0.690 ;
        RECT 14.520 0.300 14.750 0.690 ;
        RECT 0.000 -0.300 15.120 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.405 0.585 3.105 ;
        RECT 0.245 2.065 3.265 2.405 ;
        RECT 0.245 0.900 0.475 2.065 ;
        RECT 3.720 1.805 3.950 3.160 ;
        RECT 4.385 2.875 5.790 3.105 ;
        RECT 3.720 1.465 5.330 1.805 ;
        RECT 5.560 1.750 5.790 2.875 ;
        RECT 8.900 2.820 9.285 3.160 ;
        RECT 8.900 1.875 9.130 2.820 ;
        RECT 9.720 2.465 9.950 3.160 ;
        RECT 9.720 2.235 11.690 2.465 ;
        RECT 5.560 1.520 8.115 1.750 ;
        RECT 8.900 1.535 11.080 1.875 ;
        RECT 11.370 1.730 11.690 2.235 ;
        RECT 0.245 0.670 0.585 0.900 ;
        RECT 3.720 0.770 4.105 1.465 ;
        RECT 5.560 1.000 5.790 1.520 ;
        RECT 4.485 0.770 5.790 1.000 ;
        RECT 8.900 0.715 9.130 1.535 ;
        RECT 11.370 1.500 12.810 1.730 ;
        RECT 11.370 1.055 11.690 1.500 ;
        RECT 9.720 0.715 11.690 1.055 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlyc_2
MACRO gf180mcu_fd_sc_mcu7t5v0__dlyc_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlyc_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.360 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.930 1.200 3.405 1.600 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.403500 ;
    PORT
      LAYER Metal1 ;
        RECT 13.395 2.660 13.735 3.195 ;
        RECT 15.540 2.660 16.150 3.255 ;
        RECT 13.395 2.425 16.150 2.660 ;
        RECT 15.540 1.155 16.150 2.425 ;
        RECT 13.395 0.925 16.150 1.155 ;
        RECT 13.395 0.675 13.630 0.925 ;
        RECT 15.540 0.730 16.150 0.925 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 17.360 4.220 ;
        RECT 1.485 3.285 1.825 3.620 ;
        RECT 6.465 3.285 6.805 3.620 ;
        RECT 11.745 3.175 12.085 3.620 ;
        RECT 14.465 3.175 14.805 3.620 ;
        RECT 16.555 2.705 16.895 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 17.790 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 17.790 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.585 0.300 1.925 0.635 ;
        RECT 6.665 0.300 7.005 0.635 ;
        RECT 11.925 0.300 12.155 0.695 ;
        RECT 14.520 0.300 14.750 0.695 ;
        RECT 16.760 0.300 16.990 0.695 ;
        RECT 0.000 -0.300 17.360 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.405 0.585 3.105 ;
        RECT 0.245 2.065 3.265 2.405 ;
        RECT 0.245 0.900 0.475 2.065 ;
        RECT 3.720 1.805 3.950 3.160 ;
        RECT 4.385 2.875 6.260 3.105 ;
        RECT 3.720 1.465 5.800 1.805 ;
        RECT 6.030 1.750 6.260 2.875 ;
        RECT 8.900 2.820 9.285 3.160 ;
        RECT 8.900 1.875 9.130 2.820 ;
        RECT 9.720 2.465 9.950 3.160 ;
        RECT 9.720 2.235 11.690 2.465 ;
        RECT 6.030 1.520 8.115 1.750 ;
        RECT 8.900 1.535 11.080 1.875 ;
        RECT 11.370 1.760 11.690 2.235 ;
        RECT 0.245 0.670 0.585 0.900 ;
        RECT 3.720 0.770 4.105 1.465 ;
        RECT 6.030 1.000 6.260 1.520 ;
        RECT 4.485 0.770 6.260 1.000 ;
        RECT 8.900 0.715 9.130 1.535 ;
        RECT 11.370 1.530 14.690 1.760 ;
        RECT 11.370 1.055 11.690 1.530 ;
        RECT 9.720 0.715 11.690 1.055 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlyc_4
MACRO gf180mcu_fd_sc_mcu7t5v0__dlyd_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlyd_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.040 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.930 1.200 3.355 1.600 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 18.480 0.600 18.920 3.320 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 19.040 4.220 ;
        RECT 1.485 3.285 1.825 3.620 ;
        RECT 6.465 3.285 6.805 3.620 ;
        RECT 11.745 3.285 12.085 3.620 ;
        RECT 17.025 3.175 17.365 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 19.470 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 19.470 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.585 0.300 1.925 0.635 ;
        RECT 6.665 0.300 7.005 0.635 ;
        RECT 11.945 0.300 12.285 0.635 ;
        RECT 17.180 0.300 17.410 0.690 ;
        RECT 0.000 -0.300 19.040 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.405 0.585 3.105 ;
        RECT 0.245 2.065 3.265 2.405 ;
        RECT 0.245 0.900 0.475 2.065 ;
        RECT 3.720 1.805 3.950 3.160 ;
        RECT 4.385 2.875 5.790 3.105 ;
        RECT 3.720 1.465 5.330 1.805 ;
        RECT 5.560 1.750 5.790 2.875 ;
        RECT 8.900 2.820 9.285 3.160 ;
        RECT 9.665 2.875 11.070 3.105 ;
        RECT 8.900 1.805 9.130 2.820 ;
        RECT 5.560 1.520 8.115 1.750 ;
        RECT 0.245 0.670 0.585 0.900 ;
        RECT 3.720 0.770 4.105 1.465 ;
        RECT 5.560 1.000 5.790 1.520 ;
        RECT 4.485 0.770 5.790 1.000 ;
        RECT 8.900 1.465 10.610 1.805 ;
        RECT 10.840 1.750 11.070 2.875 ;
        RECT 14.180 2.820 14.565 3.160 ;
        RECT 14.180 1.875 14.410 2.820 ;
        RECT 15.000 2.465 15.230 3.160 ;
        RECT 15.000 2.235 16.880 2.465 ;
        RECT 10.840 1.520 13.395 1.750 ;
        RECT 14.180 1.535 16.360 1.875 ;
        RECT 16.650 1.625 16.880 2.235 ;
        RECT 8.900 0.715 9.130 1.465 ;
        RECT 10.840 1.000 11.070 1.520 ;
        RECT 9.765 0.770 11.070 1.000 ;
        RECT 14.180 0.715 14.410 1.535 ;
        RECT 16.650 1.395 18.185 1.625 ;
        RECT 16.650 1.000 16.880 1.395 ;
        RECT 14.945 0.770 16.880 1.000 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlyd_1
MACRO gf180mcu_fd_sc_mcu7t5v0__dlyd_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlyd_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.160 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.930 1.200 3.395 1.600 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.060800 ;
    PORT
      LAYER Metal1 ;
        RECT 18.480 0.675 18.950 3.380 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 20.160 4.220 ;
        RECT 1.485 3.285 1.825 3.620 ;
        RECT 6.465 3.285 6.805 3.620 ;
        RECT 11.745 3.285 12.085 3.620 ;
        RECT 17.460 2.530 17.690 3.620 ;
        RECT 19.500 2.530 19.730 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 20.590 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 20.590 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.585 0.300 1.925 0.635 ;
        RECT 6.665 0.300 7.005 0.635 ;
        RECT 11.945 0.300 12.285 0.635 ;
        RECT 17.180 0.300 17.410 0.690 ;
        RECT 19.600 0.300 19.830 0.690 ;
        RECT 0.000 -0.300 20.160 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.405 0.585 3.105 ;
        RECT 0.245 2.065 3.265 2.405 ;
        RECT 0.245 0.900 0.475 2.065 ;
        RECT 3.720 1.805 3.950 3.160 ;
        RECT 4.385 2.875 5.790 3.105 ;
        RECT 3.720 1.465 5.330 1.805 ;
        RECT 5.560 1.750 5.790 2.875 ;
        RECT 8.900 2.820 9.285 3.160 ;
        RECT 9.665 2.875 11.070 3.105 ;
        RECT 8.900 1.805 9.130 2.820 ;
        RECT 5.560 1.520 8.115 1.750 ;
        RECT 0.245 0.670 0.585 0.900 ;
        RECT 3.720 0.770 4.105 1.465 ;
        RECT 5.560 1.000 5.790 1.520 ;
        RECT 4.485 0.770 5.790 1.000 ;
        RECT 8.900 1.465 10.610 1.805 ;
        RECT 10.840 1.750 11.070 2.875 ;
        RECT 14.180 2.820 14.565 3.160 ;
        RECT 14.180 1.875 14.410 2.820 ;
        RECT 15.000 2.465 15.230 3.160 ;
        RECT 15.000 2.235 16.880 2.465 ;
        RECT 10.840 1.520 13.395 1.750 ;
        RECT 14.180 1.535 16.360 1.875 ;
        RECT 16.650 1.625 16.880 2.235 ;
        RECT 8.900 0.715 9.130 1.465 ;
        RECT 10.840 1.000 11.070 1.520 ;
        RECT 9.765 0.770 11.070 1.000 ;
        RECT 14.180 0.715 14.410 1.535 ;
        RECT 16.650 1.395 18.185 1.625 ;
        RECT 16.650 1.000 16.880 1.395 ;
        RECT 14.945 0.770 16.880 1.000 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlyd_2
MACRO gf180mcu_fd_sc_mcu7t5v0__dlyd_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlyd_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.400 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.930 1.200 3.355 1.600 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.121600 ;
    PORT
      LAYER Metal1 ;
        RECT 18.480 2.395 18.710 3.380 ;
        RECT 20.720 2.395 21.190 3.380 ;
        RECT 18.480 2.165 21.190 2.395 ;
        RECT 20.720 1.150 21.190 2.165 ;
        RECT 18.425 0.920 21.190 1.150 ;
        RECT 18.425 0.730 18.765 0.920 ;
        RECT 20.720 0.675 21.190 0.920 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 22.400 4.220 ;
        RECT 1.485 3.285 1.825 3.620 ;
        RECT 6.465 3.285 6.805 3.620 ;
        RECT 11.745 3.285 12.085 3.620 ;
        RECT 17.460 2.530 17.690 3.620 ;
        RECT 19.525 2.625 19.865 3.620 ;
        RECT 21.740 2.530 21.970 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 22.830 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 22.830 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.585 0.300 1.925 0.635 ;
        RECT 6.665 0.300 7.005 0.635 ;
        RECT 11.945 0.300 12.285 0.635 ;
        RECT 17.180 0.300 17.410 0.690 ;
        RECT 19.600 0.300 19.830 0.690 ;
        RECT 21.840 0.300 22.070 0.690 ;
        RECT 0.000 -0.300 22.400 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.405 0.585 3.105 ;
        RECT 0.245 2.065 3.265 2.405 ;
        RECT 0.245 0.900 0.475 2.065 ;
        RECT 3.720 1.805 3.950 3.160 ;
        RECT 4.385 2.875 5.790 3.105 ;
        RECT 3.720 1.465 5.330 1.805 ;
        RECT 5.560 1.750 5.790 2.875 ;
        RECT 8.900 2.820 9.285 3.160 ;
        RECT 9.665 2.875 11.070 3.105 ;
        RECT 8.900 1.805 9.130 2.820 ;
        RECT 5.560 1.520 8.115 1.750 ;
        RECT 0.245 0.670 0.585 0.900 ;
        RECT 3.720 0.770 4.105 1.465 ;
        RECT 5.560 1.000 5.790 1.520 ;
        RECT 4.485 0.770 5.790 1.000 ;
        RECT 8.900 1.465 10.610 1.805 ;
        RECT 10.840 1.750 11.070 2.875 ;
        RECT 14.180 2.820 14.565 3.160 ;
        RECT 14.180 1.875 14.410 2.820 ;
        RECT 15.000 2.465 15.230 3.160 ;
        RECT 15.000 2.235 16.880 2.465 ;
        RECT 10.840 1.520 13.395 1.750 ;
        RECT 14.180 1.535 16.360 1.875 ;
        RECT 16.650 1.820 16.880 2.235 ;
        RECT 16.650 1.590 20.065 1.820 ;
        RECT 8.900 0.715 9.130 1.465 ;
        RECT 10.840 1.000 11.070 1.520 ;
        RECT 9.765 0.770 11.070 1.000 ;
        RECT 14.180 0.715 14.410 1.535 ;
        RECT 16.650 1.000 16.880 1.590 ;
        RECT 14.945 0.770 16.880 1.000 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlyd_4
MACRO gf180mcu_fd_sc_mcu7t5v0__endcap
  CLASS ENDCAP PRE ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__endcap ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.120 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 1.550 4.350 ;
      LAYER Metal1 ;
        RECT 0.000 3.620 1.120 4.220 ;
        RECT 0.370 1.920 0.710 3.620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 1.550 1.760 ;
      LAYER Metal1 ;
        RECT 0.370 0.300 0.710 1.190 ;
        RECT 0.000 -0.300 1.120 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__endcap
MACRO gf180mcu_fd_sc_mcu7t5v0__fill_1
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fill_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.560 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 0.560 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 0.990 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 0.990 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.300 0.560 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__fill_1
MACRO gf180mcu_fd_sc_mcu7t5v0__fill_2
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fill_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.120 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 1.120 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 1.550 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 1.550 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.300 1.120 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__fill_2
MACRO gf180mcu_fd_sc_mcu7t5v0__fill_4
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fill_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 2.240 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 2.670 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.300 2.240 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__fill_4
MACRO gf180mcu_fd_sc_mcu7t5v0__fill_8
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fill_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 4.480 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 4.910 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.300 4.480 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__fill_8
MACRO gf180mcu_fd_sc_mcu7t5v0__fill_16
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fill_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.960 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 8.960 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 9.390 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.390 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.300 8.960 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__fill_16
MACRO gf180mcu_fd_sc_mcu7t5v0__fill_32
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fill_32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 17.920 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 18.350 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.300 17.920 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__fill_32
MACRO gf180mcu_fd_sc_mcu7t5v0__fill_64
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fill_64 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.840 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 35.840 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 36.270 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 36.270 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.300 35.840 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__fill_64
MACRO gf180mcu_fd_sc_mcu7t5v0__fillcap_4
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fillcap_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 2.240 4.220 ;
        RECT 1.765 2.490 1.995 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 2.670 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.095 ;
        RECT 0.000 -0.300 2.240 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.555 0.475 3.390 ;
        RECT 0.730 1.960 1.995 2.190 ;
        RECT 0.245 1.325 1.520 1.555 ;
        RECT 1.765 0.530 1.995 1.960 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__fillcap_4
MACRO gf180mcu_fd_sc_mcu7t5v0__fillcap_8
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fillcap_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 4.480 4.220 ;
        RECT 1.765 2.490 1.995 3.620 ;
        RECT 4.005 2.490 4.235 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 4.910 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.085 ;
        RECT 2.485 0.300 2.715 1.085 ;
        RECT 0.000 -0.300 4.480 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.555 0.475 3.390 ;
        RECT 0.730 1.960 1.995 2.190 ;
        RECT 0.245 1.325 1.520 1.555 ;
        RECT 1.765 0.530 1.995 1.960 ;
        RECT 2.485 1.555 2.715 3.390 ;
        RECT 2.970 1.960 4.235 2.190 ;
        RECT 2.485 1.325 3.760 1.555 ;
        RECT 4.005 0.530 4.235 1.960 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__fillcap_8
MACRO gf180mcu_fd_sc_mcu7t5v0__fillcap_16
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fillcap_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.960 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 8.960 4.220 ;
        RECT 1.765 2.490 1.995 3.620 ;
        RECT 4.005 2.490 4.235 3.620 ;
        RECT 6.245 2.490 6.475 3.620 ;
        RECT 8.485 2.490 8.715 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 9.390 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.390 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.070 ;
        RECT 2.485 0.300 2.715 1.070 ;
        RECT 4.725 0.300 4.955 1.070 ;
        RECT 6.965 0.300 7.195 1.070 ;
        RECT 0.000 -0.300 8.960 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.555 0.475 3.390 ;
        RECT 0.730 1.960 1.995 2.190 ;
        RECT 0.245 1.325 1.520 1.555 ;
        RECT 1.765 0.530 1.995 1.960 ;
        RECT 2.485 1.555 2.715 3.390 ;
        RECT 2.970 1.960 4.235 2.190 ;
        RECT 2.485 1.325 3.760 1.555 ;
        RECT 4.005 0.530 4.235 1.960 ;
        RECT 4.725 1.555 4.955 3.390 ;
        RECT 5.210 1.960 6.475 2.190 ;
        RECT 4.725 1.325 6.000 1.555 ;
        RECT 6.245 0.530 6.475 1.960 ;
        RECT 6.965 1.555 7.195 3.390 ;
        RECT 7.450 1.960 8.715 2.190 ;
        RECT 6.965 1.325 8.240 1.555 ;
        RECT 8.485 0.530 8.715 1.960 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__fillcap_16
MACRO gf180mcu_fd_sc_mcu7t5v0__fillcap_32
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fillcap_32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 17.920 4.220 ;
        RECT 1.765 2.490 1.995 3.620 ;
        RECT 4.005 2.490 4.235 3.620 ;
        RECT 6.245 2.490 6.475 3.620 ;
        RECT 8.485 2.490 8.715 3.620 ;
        RECT 10.725 2.490 10.955 3.620 ;
        RECT 12.965 2.490 13.195 3.620 ;
        RECT 15.205 2.490 15.435 3.620 ;
        RECT 17.445 2.490 17.675 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 18.350 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.045 ;
        RECT 2.485 0.300 2.715 1.045 ;
        RECT 4.725 0.300 4.955 1.045 ;
        RECT 6.965 0.300 7.195 1.045 ;
        RECT 9.205 0.300 9.435 1.045 ;
        RECT 11.445 0.300 11.675 1.045 ;
        RECT 13.685 0.300 13.915 1.045 ;
        RECT 15.925 0.300 16.155 1.045 ;
        RECT 0.000 -0.300 17.920 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.555 0.475 3.390 ;
        RECT 0.730 1.960 1.995 2.190 ;
        RECT 0.245 1.325 1.520 1.555 ;
        RECT 1.765 0.530 1.995 1.960 ;
        RECT 2.485 1.555 2.715 3.390 ;
        RECT 2.970 1.960 4.235 2.190 ;
        RECT 2.485 1.325 3.760 1.555 ;
        RECT 4.005 0.530 4.235 1.960 ;
        RECT 4.725 1.555 4.955 3.390 ;
        RECT 5.210 1.960 6.475 2.190 ;
        RECT 4.725 1.325 6.000 1.555 ;
        RECT 6.245 0.530 6.475 1.960 ;
        RECT 6.965 1.555 7.195 3.390 ;
        RECT 7.450 1.960 8.715 2.190 ;
        RECT 6.965 1.325 8.240 1.555 ;
        RECT 8.485 0.530 8.715 1.960 ;
        RECT 9.205 1.555 9.435 3.390 ;
        RECT 9.690 1.960 10.955 2.190 ;
        RECT 9.205 1.325 10.480 1.555 ;
        RECT 10.725 0.530 10.955 1.960 ;
        RECT 11.445 1.555 11.675 3.390 ;
        RECT 11.930 1.960 13.195 2.190 ;
        RECT 11.445 1.325 12.720 1.555 ;
        RECT 12.965 0.530 13.195 1.960 ;
        RECT 13.685 1.555 13.915 3.390 ;
        RECT 14.170 1.960 15.435 2.190 ;
        RECT 13.685 1.325 14.960 1.555 ;
        RECT 15.205 0.530 15.435 1.960 ;
        RECT 15.925 1.555 16.155 3.390 ;
        RECT 16.410 1.960 17.675 2.190 ;
        RECT 15.925 1.325 17.200 1.555 ;
        RECT 17.445 0.530 17.675 1.960 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__fillcap_32
MACRO gf180mcu_fd_sc_mcu7t5v0__fillcap_64
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fillcap_64 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.840 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 35.840 4.220 ;
        RECT 1.765 2.490 1.995 3.620 ;
        RECT 4.005 2.490 4.235 3.620 ;
        RECT 6.245 2.490 6.475 3.620 ;
        RECT 8.485 2.490 8.715 3.620 ;
        RECT 10.725 2.490 10.955 3.620 ;
        RECT 12.965 2.490 13.195 3.620 ;
        RECT 15.205 2.490 15.435 3.620 ;
        RECT 17.445 2.490 17.675 3.620 ;
        RECT 19.685 2.490 19.915 3.620 ;
        RECT 21.925 2.490 22.155 3.620 ;
        RECT 24.165 2.490 24.395 3.620 ;
        RECT 26.405 2.490 26.635 3.620 ;
        RECT 28.645 2.490 28.875 3.620 ;
        RECT 30.885 2.490 31.115 3.620 ;
        RECT 33.125 2.490 33.355 3.620 ;
        RECT 35.365 2.490 35.595 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 36.270 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 36.270 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.055 ;
        RECT 2.485 0.300 2.715 1.055 ;
        RECT 4.725 0.300 4.955 1.055 ;
        RECT 6.965 0.300 7.195 1.055 ;
        RECT 9.205 0.300 9.435 1.055 ;
        RECT 11.445 0.300 11.675 1.055 ;
        RECT 13.685 0.300 13.915 1.055 ;
        RECT 15.925 0.300 16.155 1.055 ;
        RECT 18.165 0.300 18.395 1.055 ;
        RECT 20.405 0.300 20.635 1.055 ;
        RECT 22.645 0.300 22.875 1.055 ;
        RECT 24.885 0.300 25.115 1.055 ;
        RECT 27.125 0.300 27.355 1.055 ;
        RECT 29.365 0.300 29.595 1.055 ;
        RECT 31.605 0.300 31.835 1.055 ;
        RECT 33.845 0.300 34.075 1.055 ;
        RECT 0.000 -0.300 35.840 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.555 0.475 3.390 ;
        RECT 0.730 1.960 1.995 2.190 ;
        RECT 0.245 1.325 1.520 1.555 ;
        RECT 1.765 0.530 1.995 1.960 ;
        RECT 2.485 1.555 2.715 3.390 ;
        RECT 2.970 1.960 4.235 2.190 ;
        RECT 2.485 1.325 3.760 1.555 ;
        RECT 4.005 0.530 4.235 1.960 ;
        RECT 4.725 1.555 4.955 3.390 ;
        RECT 5.210 1.960 6.475 2.190 ;
        RECT 4.725 1.325 6.000 1.555 ;
        RECT 6.245 0.530 6.475 1.960 ;
        RECT 6.965 1.555 7.195 3.390 ;
        RECT 7.450 1.960 8.715 2.190 ;
        RECT 6.965 1.325 8.240 1.555 ;
        RECT 8.485 0.530 8.715 1.960 ;
        RECT 9.205 1.555 9.435 3.390 ;
        RECT 9.690 1.960 10.955 2.190 ;
        RECT 9.205 1.325 10.480 1.555 ;
        RECT 10.725 0.530 10.955 1.960 ;
        RECT 11.445 1.555 11.675 3.390 ;
        RECT 11.930 1.960 13.195 2.190 ;
        RECT 11.445 1.325 12.720 1.555 ;
        RECT 12.965 0.530 13.195 1.960 ;
        RECT 13.685 1.555 13.915 3.390 ;
        RECT 14.170 1.960 15.435 2.190 ;
        RECT 13.685 1.325 14.960 1.555 ;
        RECT 15.205 0.530 15.435 1.960 ;
        RECT 15.925 1.555 16.155 3.390 ;
        RECT 16.410 1.960 17.675 2.190 ;
        RECT 15.925 1.325 17.200 1.555 ;
        RECT 17.445 0.530 17.675 1.960 ;
        RECT 18.165 1.555 18.395 3.390 ;
        RECT 18.650 1.960 19.915 2.190 ;
        RECT 18.165 1.325 19.440 1.555 ;
        RECT 19.685 0.530 19.915 1.960 ;
        RECT 20.405 1.555 20.635 3.390 ;
        RECT 20.890 1.960 22.155 2.190 ;
        RECT 20.405 1.325 21.680 1.555 ;
        RECT 21.925 0.530 22.155 1.960 ;
        RECT 22.645 1.555 22.875 3.390 ;
        RECT 23.130 1.960 24.395 2.190 ;
        RECT 22.645 1.325 23.920 1.555 ;
        RECT 24.165 0.530 24.395 1.960 ;
        RECT 24.885 1.555 25.115 3.390 ;
        RECT 25.370 1.960 26.635 2.190 ;
        RECT 24.885 1.325 26.160 1.555 ;
        RECT 26.405 0.530 26.635 1.960 ;
        RECT 27.125 1.555 27.355 3.390 ;
        RECT 27.610 1.960 28.875 2.190 ;
        RECT 27.125 1.325 28.400 1.555 ;
        RECT 28.645 0.530 28.875 1.960 ;
        RECT 29.365 1.555 29.595 3.390 ;
        RECT 29.850 1.960 31.115 2.190 ;
        RECT 29.365 1.325 30.640 1.555 ;
        RECT 30.885 0.530 31.115 1.960 ;
        RECT 31.605 1.555 31.835 3.390 ;
        RECT 32.090 1.960 33.355 2.190 ;
        RECT 31.605 1.325 32.880 1.555 ;
        RECT 33.125 0.530 33.355 1.960 ;
        RECT 33.845 1.555 34.075 3.390 ;
        RECT 34.330 1.960 35.595 2.190 ;
        RECT 33.845 1.325 35.120 1.555 ;
        RECT 35.365 0.530 35.595 1.960 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__fillcap_64
MACRO gf180mcu_fd_sc_mcu7t5v0__filltie
  CLASS core WELLTAP ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__filltie ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.120 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 1.550 4.350 ;
      LAYER Metal1 ;
        RECT 0.000 3.620 1.120 4.220 ;
        RECT 0.390 1.930 0.730 3.620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 1.550 1.760 ;
      LAYER Metal1 ;
        RECT 0.390 0.300 0.730 1.185 ;
        RECT 0.000 -0.300 1.120 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__filltie
MACRO gf180mcu_fd_sc_mcu7t5v0__hold
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__hold ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.040 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN Z
    DIRECTION INOUT ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.451200 ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 1.560 0.575 2.895 ;
        RECT 0.245 1.155 3.950 1.560 ;
        RECT 0.245 0.565 0.475 1.155 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.040 4.220 ;
        RECT 3.225 2.535 3.455 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 5.470 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 5.470 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.225 0.300 3.455 0.925 ;
        RECT 0.000 -0.300 5.040 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 4.245 2.185 4.575 3.180 ;
        RECT 2.450 1.885 4.575 2.185 ;
        RECT 4.345 0.575 4.575 1.885 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__hold
MACRO gf180mcu_fd_sc_mcu7t5v0__icgtn_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__icgtn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.360 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.394000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.025 1.680 14.255 2.195 ;
        RECT 13.570 1.590 14.255 1.680 ;
        RECT 11.810 1.450 14.255 1.590 ;
        RECT 11.810 1.210 13.865 1.450 ;
    END
  END CLKN
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.699500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.320 2.150 2.730 3.370 ;
        RECT 1.845 1.770 2.730 2.150 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.699500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.270 1.770 1.570 2.150 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.811800 ;
    PORT
      LAYER Metal1 ;
        RECT 16.300 0.630 17.035 3.270 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 17.360 4.220 ;
        RECT 0.345 2.480 0.575 3.620 ;
        RECT 6.300 2.790 6.530 3.620 ;
        RECT 9.110 2.470 9.340 3.620 ;
        RECT 12.800 2.460 13.030 3.620 ;
        RECT 15.345 2.425 15.685 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.775 17.790 4.350 ;
        RECT -0.430 1.760 4.735 1.775 ;
        RECT 10.880 1.760 17.790 1.775 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 4.735 1.760 10.880 1.775 ;
        RECT -0.430 -0.430 17.790 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 1.060 ;
        RECT 6.065 0.300 6.405 1.075 ;
        RECT 9.105 0.300 9.445 1.075 ;
        RECT 12.665 0.300 13.005 0.760 ;
        RECT 14.905 0.300 15.245 0.760 ;
        RECT 15.680 0.300 15.910 1.095 ;
        RECT 0.000 -0.300 17.360 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 6.810 3.160 8.790 3.390 ;
        RECT 3.810 2.560 4.040 3.125 ;
        RECT 6.810 2.560 7.040 3.160 ;
        RECT 3.000 2.330 7.040 2.560 ;
        RECT 0.190 1.290 2.115 1.520 ;
        RECT 0.190 0.845 0.530 1.290 ;
        RECT 1.885 1.075 2.115 1.290 ;
        RECT 3.000 1.075 3.230 2.330 ;
        RECT 7.320 2.100 7.550 2.900 ;
        RECT 3.460 1.870 7.550 2.100 ;
        RECT 3.460 1.420 3.690 1.870 ;
        RECT 1.885 0.845 2.770 1.075 ;
        RECT 3.000 0.845 3.890 1.075 ;
        RECT 7.320 0.780 7.550 1.870 ;
        RECT 8.040 1.575 8.270 2.900 ;
        RECT 8.560 1.820 8.790 3.160 ;
        RECT 10.180 3.160 12.570 3.390 ;
        RECT 8.040 1.340 9.910 1.575 ;
        RECT 8.040 0.780 8.270 1.340 ;
        RECT 10.180 0.780 10.510 3.160 ;
        RECT 11.780 2.495 12.010 2.930 ;
        RECT 10.860 2.260 12.010 2.495 ;
        RECT 10.860 0.760 11.090 2.260 ;
        RECT 12.340 2.140 12.570 3.160 ;
        RECT 12.340 1.910 13.630 2.140 ;
        RECT 14.560 2.130 14.790 3.180 ;
        RECT 14.560 1.790 16.070 2.130 ;
        RECT 14.560 1.220 14.790 1.790 ;
        RECT 14.340 0.990 14.790 1.220 ;
        RECT 14.340 0.760 14.570 0.990 ;
        RECT 10.860 0.530 11.975 0.760 ;
        RECT 13.785 0.530 14.570 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__icgtn_1
MACRO gf180mcu_fd_sc_mcu7t5v0__icgtn_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__icgtn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.480 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.725000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.985 1.590 14.215 2.250 ;
        RECT 11.810 1.210 14.215 1.590 ;
    END
  END CLKN
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.699500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.340 2.150 2.750 3.370 ;
        RECT 1.865 1.770 2.750 2.150 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.699500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.290 1.770 1.590 2.150 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.962000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.455 2.710 16.795 3.305 ;
        RECT 16.455 2.370 17.830 2.710 ;
        RECT 17.450 1.415 17.830 2.370 ;
        RECT 16.750 1.145 17.830 1.415 ;
        RECT 16.750 0.600 17.220 1.145 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 18.480 4.220 ;
        RECT 0.345 2.480 0.575 3.620 ;
        RECT 6.300 2.790 6.530 3.620 ;
        RECT 9.110 2.470 9.340 3.620 ;
        RECT 12.800 2.695 13.030 3.620 ;
        RECT 15.490 2.610 15.720 3.620 ;
        RECT 17.530 3.020 17.760 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.775 18.910 4.350 ;
        RECT -0.430 1.760 4.760 1.775 ;
        RECT 10.710 1.760 18.910 1.775 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 4.760 1.760 10.710 1.775 ;
        RECT -0.430 -0.430 18.910 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 1.060 ;
        RECT 6.065 0.300 6.405 1.075 ;
        RECT 9.105 0.300 9.445 1.075 ;
        RECT 12.665 0.300 13.005 0.760 ;
        RECT 14.905 0.300 15.245 0.760 ;
        RECT 15.680 0.300 15.910 1.090 ;
        RECT 17.920 0.300 18.150 0.915 ;
        RECT 0.000 -0.300 18.480 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.810 2.560 4.040 3.265 ;
        RECT 6.810 3.160 8.790 3.390 ;
        RECT 6.810 2.560 7.040 3.160 ;
        RECT 3.000 2.330 7.040 2.560 ;
        RECT 0.190 1.290 2.115 1.520 ;
        RECT 0.190 0.845 0.530 1.290 ;
        RECT 1.885 1.075 2.115 1.290 ;
        RECT 3.000 1.075 3.230 2.330 ;
        RECT 7.320 2.100 7.550 2.900 ;
        RECT 3.460 1.870 7.550 2.100 ;
        RECT 3.460 1.420 3.690 1.870 ;
        RECT 1.885 0.845 2.770 1.075 ;
        RECT 3.000 0.845 3.890 1.075 ;
        RECT 7.320 0.780 7.550 1.870 ;
        RECT 8.040 1.575 8.270 2.900 ;
        RECT 8.560 1.820 8.790 3.160 ;
        RECT 10.180 3.160 12.570 3.390 ;
        RECT 8.040 1.340 9.910 1.575 ;
        RECT 8.040 0.780 8.270 1.340 ;
        RECT 10.180 0.780 10.510 3.160 ;
        RECT 11.780 2.495 12.010 2.930 ;
        RECT 10.860 2.260 12.010 2.495 ;
        RECT 10.860 0.760 11.090 2.260 ;
        RECT 12.340 2.140 12.570 3.160 ;
        RECT 14.560 2.140 14.790 3.180 ;
        RECT 12.340 1.910 13.630 2.140 ;
        RECT 14.560 2.130 17.190 2.140 ;
        RECT 14.445 1.790 17.190 2.130 ;
        RECT 14.445 0.990 14.790 1.790 ;
        RECT 14.445 0.760 14.675 0.990 ;
        RECT 10.860 0.530 11.885 0.760 ;
        RECT 13.785 0.530 14.675 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__icgtn_2
MACRO gf180mcu_fd_sc_mcu7t5v0__icgtn_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__icgtn_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.720 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.725000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.025 1.680 14.255 2.195 ;
        RECT 13.570 1.590 14.255 1.680 ;
        RECT 11.810 1.450 14.255 1.590 ;
        RECT 11.810 1.210 13.865 1.450 ;
    END
  END CLKN
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.699500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.340 2.120 2.750 3.370 ;
        RECT 1.865 1.800 2.750 2.120 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.699500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.290 1.800 1.590 2.120 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.924000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.510 2.710 16.740 3.180 ;
        RECT 18.550 2.710 18.780 3.180 ;
        RECT 16.510 2.370 20.070 2.710 ;
        RECT 19.690 1.535 20.070 2.370 ;
        RECT 16.750 1.265 20.070 1.535 ;
        RECT 16.750 0.600 17.220 1.265 ;
        RECT 19.040 0.600 19.470 1.265 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 20.720 4.220 ;
        RECT 0.345 2.480 0.575 3.620 ;
        RECT 6.300 2.790 6.530 3.620 ;
        RECT 9.110 2.470 9.340 3.620 ;
        RECT 12.800 2.645 13.030 3.620 ;
        RECT 15.490 2.645 15.720 3.620 ;
        RECT 17.530 3.020 17.760 3.620 ;
        RECT 19.570 3.020 19.800 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.775 21.150 4.350 ;
        RECT -0.430 1.760 4.760 1.775 ;
        RECT 10.710 1.760 21.150 1.775 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 4.760 1.760 10.710 1.775 ;
        RECT -0.430 -0.430 21.150 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 1.060 ;
        RECT 6.065 0.300 6.405 1.075 ;
        RECT 9.105 0.300 9.445 1.075 ;
        RECT 12.665 0.300 13.005 0.760 ;
        RECT 14.905 0.300 15.245 0.760 ;
        RECT 15.680 0.300 15.910 1.090 ;
        RECT 17.920 0.300 18.150 0.975 ;
        RECT 20.160 0.300 20.390 0.975 ;
        RECT 0.000 -0.300 20.720 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.810 2.560 4.040 3.265 ;
        RECT 6.810 3.160 8.790 3.390 ;
        RECT 6.810 2.560 7.040 3.160 ;
        RECT 3.000 2.330 7.040 2.560 ;
        RECT 0.190 1.305 2.115 1.540 ;
        RECT 0.190 0.845 0.530 1.305 ;
        RECT 1.885 1.075 2.115 1.305 ;
        RECT 3.000 1.075 3.230 2.330 ;
        RECT 7.320 2.100 7.550 2.900 ;
        RECT 3.460 1.870 7.550 2.100 ;
        RECT 3.460 1.420 3.690 1.870 ;
        RECT 1.885 0.845 2.770 1.075 ;
        RECT 3.000 0.845 3.890 1.075 ;
        RECT 7.320 0.780 7.550 1.870 ;
        RECT 8.040 1.575 8.270 2.900 ;
        RECT 8.560 1.820 8.790 3.160 ;
        RECT 10.180 3.160 12.570 3.390 ;
        RECT 8.040 1.340 9.910 1.575 ;
        RECT 8.040 0.780 8.270 1.340 ;
        RECT 10.180 0.780 10.510 3.160 ;
        RECT 11.780 2.495 12.010 2.930 ;
        RECT 10.860 2.260 12.010 2.495 ;
        RECT 10.860 0.760 11.090 2.260 ;
        RECT 12.340 2.140 12.570 3.160 ;
        RECT 14.560 2.140 14.790 3.180 ;
        RECT 12.340 1.910 13.630 2.140 ;
        RECT 14.560 1.790 19.280 2.140 ;
        RECT 14.560 1.220 14.790 1.790 ;
        RECT 14.340 0.990 14.790 1.220 ;
        RECT 14.340 0.760 14.570 0.990 ;
        RECT 10.860 0.530 11.975 0.760 ;
        RECT 13.785 0.530 14.570 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__icgtn_4
MACRO gf180mcu_fd_sc_mcu7t5v0__icgtp_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__icgtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.680 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.388000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.215 1.590 11.065 1.765 ;
        RECT 10.215 1.535 12.755 1.590 ;
        RECT 10.785 1.210 12.755 1.535 ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.699500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.340 2.150 2.750 3.370 ;
        RECT 1.865 1.770 2.750 2.150 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.699500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.290 1.770 1.590 2.150 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.814000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.160 2.330 15.230 3.270 ;
        RECT 14.780 1.120 15.230 2.330 ;
        RECT 14.700 0.560 15.230 1.120 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 15.680 4.220 ;
        RECT 0.345 2.480 0.575 3.620 ;
        RECT 6.245 2.845 6.585 3.620 ;
        RECT 9.690 2.920 9.920 3.620 ;
        RECT 11.635 2.460 11.865 3.620 ;
        RECT 13.700 2.900 13.930 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.775 16.110 4.350 ;
        RECT -0.430 1.760 4.760 1.775 ;
        RECT 7.750 1.760 16.110 1.775 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 4.760 1.760 7.750 1.775 ;
        RECT -0.430 -0.430 16.110 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.995 ;
        RECT 6.065 0.300 6.405 1.075 ;
        RECT 9.820 0.300 10.050 0.845 ;
        RECT 13.700 0.300 13.930 0.805 ;
        RECT 0.000 -0.300 15.680 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 7.320 3.160 9.395 3.390 ;
        RECT 3.810 2.560 4.040 3.125 ;
        RECT 3.000 2.330 5.435 2.560 ;
        RECT 0.190 1.225 2.115 1.460 ;
        RECT 0.190 0.765 0.530 1.225 ;
        RECT 1.885 0.995 2.115 1.225 ;
        RECT 3.000 0.995 3.230 2.330 ;
        RECT 3.460 1.870 4.935 2.100 ;
        RECT 3.460 1.445 3.690 1.870 ;
        RECT 5.205 1.575 5.435 2.330 ;
        RECT 7.320 2.035 7.550 3.160 ;
        RECT 8.645 2.035 8.930 2.850 ;
        RECT 9.165 2.690 9.395 3.160 ;
        RECT 10.200 3.160 11.405 3.390 ;
        RECT 10.200 2.690 10.430 3.160 ;
        RECT 9.165 2.455 10.430 2.690 ;
        RECT 10.715 2.225 10.945 2.850 ;
        RECT 5.685 1.805 7.550 2.035 ;
        RECT 5.205 1.340 7.080 1.575 ;
        RECT 1.885 0.765 2.770 0.995 ;
        RECT 3.000 0.765 3.890 0.995 ;
        RECT 7.320 0.780 7.550 1.805 ;
        RECT 7.915 1.805 8.930 2.035 ;
        RECT 9.245 1.995 10.945 2.225 ;
        RECT 11.175 2.225 11.405 3.160 ;
        RECT 12.680 2.670 12.910 3.250 ;
        RECT 12.680 2.440 13.875 2.670 ;
        RECT 11.175 2.210 12.265 2.225 ;
        RECT 11.175 1.995 13.415 2.210 ;
        RECT 7.915 0.760 8.275 1.805 ;
        RECT 9.245 1.305 9.485 1.995 ;
        RECT 12.010 1.965 13.415 1.995 ;
        RECT 13.645 2.025 13.875 2.440 ;
        RECT 13.645 1.685 14.550 2.025 ;
        RECT 13.645 1.535 13.875 1.685 ;
        RECT 9.245 1.075 10.510 1.305 ;
        RECT 10.280 0.760 10.510 1.075 ;
        RECT 13.010 1.265 13.875 1.535 ;
        RECT 13.010 0.760 13.240 1.265 ;
        RECT 7.915 0.530 9.075 0.760 ;
        RECT 10.280 0.530 11.235 0.760 ;
        RECT 11.595 0.530 13.240 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__icgtp_1
MACRO gf180mcu_fd_sc_mcu7t5v0__icgtp_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__icgtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.800 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.679000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.110 1.590 10.970 1.765 ;
        RECT 10.110 1.535 12.755 1.590 ;
        RECT 10.740 1.210 12.755 1.535 ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.699500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.340 2.120 2.750 3.370 ;
        RECT 1.865 1.800 2.750 2.120 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.699500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.290 1.800 1.590 2.120 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.118000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.660 2.740 15.020 3.380 ;
        RECT 14.660 2.400 15.580 2.740 ;
        RECT 15.220 1.080 15.580 2.400 ;
        RECT 14.555 0.600 15.580 1.080 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 16.800 4.220 ;
        RECT 0.290 2.535 0.630 3.620 ;
        RECT 6.280 2.505 6.510 3.620 ;
        RECT 9.690 2.920 9.920 3.620 ;
        RECT 11.635 2.570 11.865 3.620 ;
        RECT 13.645 2.815 13.985 3.620 ;
        RECT 15.870 2.530 16.100 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.775 17.230 4.350 ;
        RECT -0.430 1.760 4.760 1.775 ;
        RECT 7.750 1.760 17.230 1.775 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 4.760 1.760 7.750 1.775 ;
        RECT -0.430 -0.430 17.230 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.995 ;
        RECT 6.065 0.300 6.405 1.075 ;
        RECT 9.820 0.300 10.050 0.845 ;
        RECT 13.700 0.300 13.930 0.845 ;
        RECT 15.885 0.300 16.235 0.750 ;
        RECT 0.000 -0.300 16.800 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.810 2.560 4.040 3.265 ;
        RECT 7.320 3.160 9.395 3.390 ;
        RECT 3.000 2.330 5.435 2.560 ;
        RECT 0.190 1.225 2.115 1.460 ;
        RECT 0.190 0.765 0.530 1.225 ;
        RECT 1.885 0.995 2.115 1.225 ;
        RECT 3.000 0.995 3.230 2.330 ;
        RECT 3.460 1.870 4.935 2.100 ;
        RECT 3.460 1.445 3.690 1.870 ;
        RECT 5.205 1.575 5.435 2.330 ;
        RECT 7.320 2.035 7.550 3.160 ;
        RECT 8.645 2.035 8.930 2.850 ;
        RECT 9.165 2.690 9.395 3.160 ;
        RECT 10.200 3.160 11.405 3.390 ;
        RECT 10.200 2.690 10.430 3.160 ;
        RECT 9.165 2.455 10.430 2.690 ;
        RECT 10.715 2.225 10.945 2.850 ;
        RECT 5.685 1.805 7.550 2.035 ;
        RECT 5.205 1.340 7.080 1.575 ;
        RECT 1.885 0.765 2.770 0.995 ;
        RECT 3.000 0.765 3.890 0.995 ;
        RECT 7.320 0.780 7.550 1.805 ;
        RECT 7.915 1.805 8.930 2.035 ;
        RECT 9.175 1.995 10.945 2.225 ;
        RECT 11.175 2.125 11.405 3.160 ;
        RECT 12.680 2.585 12.910 3.380 ;
        RECT 12.680 2.355 13.875 2.585 ;
        RECT 7.915 0.760 8.275 1.805 ;
        RECT 9.175 1.305 9.415 1.995 ;
        RECT 11.175 1.895 13.415 2.125 ;
        RECT 13.645 1.825 13.875 2.355 ;
        RECT 13.645 1.595 14.970 1.825 ;
        RECT 13.645 1.535 13.875 1.595 ;
        RECT 9.175 1.075 10.510 1.305 ;
        RECT 10.280 0.760 10.510 1.075 ;
        RECT 13.010 1.265 13.875 1.535 ;
        RECT 13.010 0.760 13.240 1.265 ;
        RECT 7.915 0.530 9.075 0.760 ;
        RECT 10.280 0.530 11.235 0.760 ;
        RECT 11.595 0.530 13.240 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__icgtp_2
MACRO gf180mcu_fd_sc_mcu7t5v0__icgtp_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__icgtp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.040 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.685000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.105 1.590 11.065 1.765 ;
        RECT 10.105 1.535 12.755 1.590 ;
        RECT 10.785 1.210 12.755 1.535 ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.699500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.330 2.150 2.710 3.270 ;
        RECT 1.865 1.770 2.710 2.150 ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.699500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.290 1.770 1.590 2.150 ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.924000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.700 2.710 14.975 3.195 ;
        RECT 16.760 2.710 16.990 3.195 ;
        RECT 14.700 2.330 18.390 2.710 ;
        RECT 18.010 1.535 18.390 2.330 ;
        RECT 14.820 1.265 18.390 1.535 ;
        RECT 14.820 0.705 15.050 1.265 ;
        RECT 17.060 0.705 17.290 1.265 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 19.040 4.220 ;
        RECT 0.345 2.480 0.575 3.620 ;
        RECT 6.280 2.605 6.510 3.620 ;
        RECT 9.690 2.920 9.920 3.620 ;
        RECT 11.635 2.760 11.865 3.620 ;
        RECT 13.700 3.040 13.930 3.620 ;
        RECT 15.740 3.040 15.970 3.620 ;
        RECT 17.780 3.045 18.010 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.775 19.470 4.350 ;
        RECT -0.430 1.760 4.760 1.775 ;
        RECT 7.750 1.760 19.470 1.775 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 4.760 1.760 7.750 1.775 ;
        RECT -0.430 -0.430 19.470 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.995 ;
        RECT 6.065 0.300 6.405 1.075 ;
        RECT 9.820 0.300 10.050 0.845 ;
        RECT 13.700 0.300 13.930 0.805 ;
        RECT 15.940 0.300 16.170 0.805 ;
        RECT 18.180 0.300 18.410 0.805 ;
        RECT 0.000 -0.300 19.040 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 7.320 3.160 9.395 3.390 ;
        RECT 3.810 2.560 4.040 3.125 ;
        RECT 3.000 2.330 5.435 2.560 ;
        RECT 0.190 1.225 2.115 1.460 ;
        RECT 0.190 0.765 0.530 1.225 ;
        RECT 1.885 0.995 2.115 1.225 ;
        RECT 3.000 0.995 3.230 2.330 ;
        RECT 3.460 1.870 4.935 2.100 ;
        RECT 3.460 1.445 3.690 1.870 ;
        RECT 5.205 1.575 5.435 2.330 ;
        RECT 7.320 2.035 7.550 3.160 ;
        RECT 8.645 2.035 8.930 2.850 ;
        RECT 9.165 2.690 9.395 3.160 ;
        RECT 10.200 3.160 11.405 3.390 ;
        RECT 10.200 2.690 10.430 3.160 ;
        RECT 9.165 2.455 10.430 2.690 ;
        RECT 10.715 2.225 10.945 2.850 ;
        RECT 5.685 1.805 7.550 2.035 ;
        RECT 5.205 1.340 7.080 1.575 ;
        RECT 1.885 0.765 2.770 0.995 ;
        RECT 3.000 0.765 3.890 0.995 ;
        RECT 7.320 0.780 7.550 1.805 ;
        RECT 7.915 1.805 8.930 2.035 ;
        RECT 9.175 1.995 10.945 2.225 ;
        RECT 11.175 2.225 11.405 3.160 ;
        RECT 12.680 2.685 12.910 3.265 ;
        RECT 12.680 2.455 13.930 2.685 ;
        RECT 11.175 1.995 13.415 2.225 ;
        RECT 7.915 0.760 8.275 1.805 ;
        RECT 9.175 1.305 9.415 1.995 ;
        RECT 13.075 1.965 13.415 1.995 ;
        RECT 13.700 2.095 13.930 2.455 ;
        RECT 13.700 1.825 17.570 2.095 ;
        RECT 13.700 1.535 13.930 1.825 ;
        RECT 9.175 1.075 10.510 1.305 ;
        RECT 10.280 0.760 10.510 1.075 ;
        RECT 13.105 1.265 13.930 1.535 ;
        RECT 13.105 0.760 13.335 1.265 ;
        RECT 7.915 0.530 9.075 0.760 ;
        RECT 10.280 0.530 11.235 0.760 ;
        RECT 11.595 0.530 13.335 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__icgtp_4
MACRO gf180mcu_fd_sc_mcu7t5v0__inv_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__inv_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 1.200 1.035 2.200 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 0.530 1.595 3.390 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 2.240 4.220 ;
        RECT 0.345 2.530 0.575 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 2.670 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.160 ;
        RECT 0.000 -0.300 2.240 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__inv_1
MACRO gf180mcu_fd_sc_mcu7t5v0__inv_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__inv_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 1.705 2.150 2.120 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.366000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.220 2.680 1.670 3.390 ;
        RECT 1.220 2.360 2.680 2.680 ;
        RECT 2.380 1.475 2.680 2.360 ;
        RECT 1.395 1.220 2.680 1.475 ;
        RECT 1.395 0.530 1.625 1.220 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 3.360 4.220 ;
        RECT 0.245 2.640 0.475 3.620 ;
        RECT 2.515 2.930 2.745 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 3.790 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 3.790 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 0.950 ;
        RECT 2.515 0.300 2.745 0.950 ;
        RECT 0.000 -0.300 3.360 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__inv_2
MACRO gf180mcu_fd_sc_mcu7t5v0__inv_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__inv_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.306000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.410 1.760 3.015 2.120 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.202400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 2.680 1.595 3.390 ;
        RECT 3.410 2.680 3.835 3.390 ;
        RECT 1.365 2.360 3.835 2.680 ;
        RECT 3.410 1.525 3.835 2.360 ;
        RECT 1.365 1.290 3.835 1.525 ;
        RECT 1.365 0.530 1.595 1.290 ;
        RECT 3.410 0.530 3.835 1.290 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 4.480 4.220 ;
        RECT 0.245 2.530 0.475 3.620 ;
        RECT 2.485 2.985 2.715 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 4.910 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.160 ;
        RECT 2.485 0.300 2.715 1.055 ;
        RECT 0.000 -0.300 4.480 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__inv_3
MACRO gf180mcu_fd_sc_mcu7t5v0__inv_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__inv_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.408000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.370 1.740 1.950 2.150 ;
        RECT 3.035 1.740 4.315 2.150 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.609600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 2.770 1.595 3.390 ;
        RECT 3.605 2.770 3.835 3.390 ;
        RECT 1.365 2.390 3.835 2.770 ;
        RECT 2.330 1.440 2.710 2.390 ;
        RECT 1.365 1.060 3.835 1.440 ;
        RECT 1.365 0.675 1.595 1.060 ;
        RECT 3.605 0.675 3.835 1.060 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.600 4.220 ;
        RECT 0.245 2.615 0.475 3.620 ;
        RECT 2.485 3.130 2.715 3.620 ;
        RECT 4.725 2.620 4.955 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 6.030 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 0.970 ;
        RECT 2.485 0.300 2.715 0.775 ;
        RECT 4.725 0.300 4.955 0.975 ;
        RECT 0.000 -0.300 5.600 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__inv_4
MACRO gf180mcu_fd_sc_mcu7t5v0__inv_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__inv_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 8.816000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 1.765 4.260 2.120 ;
        RECT 5.320 1.765 8.960 2.120 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.219200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 2.675 1.595 3.380 ;
        RECT 3.605 2.675 3.835 3.380 ;
        RECT 5.845 2.680 6.075 3.380 ;
        RECT 8.085 2.680 8.315 3.380 ;
        RECT 5.845 2.675 8.315 2.680 ;
        RECT 1.365 2.375 8.315 2.675 ;
        RECT 4.570 1.535 4.950 2.375 ;
        RECT 1.365 1.235 8.315 1.535 ;
        RECT 1.365 0.675 1.595 1.235 ;
        RECT 3.605 0.675 3.835 1.235 ;
        RECT 5.845 0.675 6.075 1.235 ;
        RECT 8.085 0.675 8.315 1.235 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 10.080 4.220 ;
        RECT 0.245 2.655 0.475 3.620 ;
        RECT 2.485 2.950 2.715 3.620 ;
        RECT 4.725 2.950 4.955 3.620 ;
        RECT 6.965 2.950 7.195 3.620 ;
        RECT 9.205 2.650 9.435 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 10.510 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.015 ;
        RECT 2.485 0.300 2.715 0.995 ;
        RECT 4.725 0.300 4.955 0.995 ;
        RECT 6.965 0.300 7.195 0.995 ;
        RECT 9.205 0.300 9.435 1.015 ;
        RECT 0.000 -0.300 10.080 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__inv_8
MACRO gf180mcu_fd_sc_mcu7t5v0__inv_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__inv_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 13.224000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.640 1.765 6.155 2.150 ;
        RECT 7.800 1.765 13.310 2.150 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.096800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 2.960 1.595 3.390 ;
        RECT 3.505 2.960 3.735 3.390 ;
        RECT 5.745 2.960 5.975 3.390 ;
        RECT 7.985 2.960 8.215 3.390 ;
        RECT 10.225 2.960 10.455 3.390 ;
        RECT 12.465 2.960 12.695 3.390 ;
        RECT 1.365 2.535 12.695 2.960 ;
        RECT 1.365 2.520 7.450 2.535 ;
        RECT 6.550 1.450 7.450 2.520 ;
        RECT 1.365 1.010 12.795 1.450 ;
        RECT 1.365 0.675 1.595 1.010 ;
        RECT 3.605 0.675 3.835 1.010 ;
        RECT 5.845 0.675 6.075 1.010 ;
        RECT 8.085 0.675 8.315 1.010 ;
        RECT 10.325 0.675 10.555 1.010 ;
        RECT 12.565 0.675 12.795 1.010 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 14.560 4.220 ;
        RECT 0.245 2.680 0.475 3.620 ;
        RECT 2.385 3.210 2.615 3.620 ;
        RECT 4.625 3.210 4.855 3.620 ;
        RECT 6.865 3.210 7.095 3.620 ;
        RECT 9.105 3.210 9.335 3.620 ;
        RECT 11.345 3.210 11.575 3.620 ;
        RECT 13.585 2.680 13.815 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 14.990 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.015 ;
        RECT 2.485 0.300 2.715 0.690 ;
        RECT 4.725 0.300 4.955 0.690 ;
        RECT 6.965 0.300 7.195 0.690 ;
        RECT 9.205 0.300 9.435 0.690 ;
        RECT 11.445 0.300 11.675 0.690 ;
        RECT 13.685 0.300 13.915 1.015 ;
        RECT 0.000 -0.300 14.560 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__inv_12
MACRO gf180mcu_fd_sc_mcu7t5v0__inv_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__inv_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.040 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 17.632000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.620 1.765 8.510 2.190 ;
        RECT 10.015 1.765 17.920 2.190 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.462399 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.000 1.595 3.390 ;
        RECT 3.505 3.000 3.735 3.390 ;
        RECT 5.745 3.000 5.975 3.390 ;
        RECT 8.080 3.000 8.310 3.390 ;
        RECT 10.225 3.000 10.455 3.390 ;
        RECT 12.465 3.000 12.695 3.390 ;
        RECT 14.705 3.000 14.935 3.390 ;
        RECT 16.945 3.000 17.175 3.390 ;
        RECT 1.365 2.420 17.175 3.000 ;
        RECT 8.790 1.445 9.690 2.420 ;
        RECT 1.365 0.865 17.275 1.445 ;
        RECT 1.365 0.675 1.625 0.865 ;
        RECT 3.605 0.675 3.835 0.865 ;
        RECT 5.845 0.675 6.075 0.865 ;
        RECT 8.085 0.675 8.315 0.865 ;
        RECT 10.325 0.675 10.555 0.865 ;
        RECT 12.565 0.675 12.795 0.865 ;
        RECT 14.805 0.675 15.035 0.865 ;
        RECT 17.045 0.675 17.275 0.865 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 19.040 4.220 ;
        RECT 0.245 2.680 0.475 3.620 ;
        RECT 2.385 3.230 2.615 3.620 ;
        RECT 4.625 3.230 4.855 3.620 ;
        RECT 6.865 3.230 7.095 3.620 ;
        RECT 9.105 3.230 9.335 3.620 ;
        RECT 11.345 3.230 11.575 3.620 ;
        RECT 13.585 3.230 13.815 3.620 ;
        RECT 15.825 3.230 16.055 3.620 ;
        RECT 18.065 2.680 18.295 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 19.470 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 19.470 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.015 ;
        RECT 2.430 0.300 2.770 0.635 ;
        RECT 4.670 0.300 5.010 0.635 ;
        RECT 6.910 0.300 7.250 0.635 ;
        RECT 9.150 0.300 9.490 0.635 ;
        RECT 11.390 0.300 11.730 0.635 ;
        RECT 13.630 0.300 13.970 0.635 ;
        RECT 15.870 0.300 16.210 0.635 ;
        RECT 18.165 0.300 18.395 1.015 ;
        RECT 0.000 -0.300 19.040 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__inv_16
MACRO gf180mcu_fd_sc_mcu7t5v0__inv_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__inv_20 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.520 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 22.039999 ;
    PORT
      LAYER Metal1 ;
        RECT 0.610 1.765 8.020 2.150 ;
        RECT 14.985 1.765 22.375 2.150 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 11.828000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 3.055 1.595 3.375 ;
        RECT 3.505 3.055 3.735 3.375 ;
        RECT 5.745 3.055 5.975 3.375 ;
        RECT 7.985 3.055 8.215 3.375 ;
        RECT 10.225 3.055 10.455 3.375 ;
        RECT 12.465 3.055 12.695 3.375 ;
        RECT 14.705 3.055 14.935 3.375 ;
        RECT 16.945 3.055 17.175 3.375 ;
        RECT 19.185 3.055 19.415 3.375 ;
        RECT 21.425 3.055 21.655 3.375 ;
        RECT 1.365 2.380 21.655 3.055 ;
        RECT 8.395 2.315 14.665 2.380 ;
        RECT 11.030 1.605 11.930 2.315 ;
        RECT 8.415 1.535 14.770 1.605 ;
        RECT 1.310 0.865 21.755 1.535 ;
        RECT 1.310 0.730 1.650 0.865 ;
        RECT 3.605 0.675 3.835 0.865 ;
        RECT 5.845 0.675 6.075 0.865 ;
        RECT 8.085 0.675 8.315 0.865 ;
        RECT 10.325 0.675 10.555 0.865 ;
        RECT 12.565 0.675 12.795 0.865 ;
        RECT 14.805 0.675 15.035 0.865 ;
        RECT 17.045 0.675 17.275 0.865 ;
        RECT 19.285 0.675 19.515 0.865 ;
        RECT 21.525 0.675 21.755 0.865 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 23.520 4.220 ;
        RECT 0.245 2.640 0.475 3.620 ;
        RECT 2.330 3.285 2.670 3.620 ;
        RECT 4.570 3.285 4.910 3.620 ;
        RECT 6.810 3.285 7.150 3.620 ;
        RECT 9.050 3.285 9.390 3.620 ;
        RECT 11.290 3.285 11.630 3.620 ;
        RECT 13.530 3.285 13.870 3.620 ;
        RECT 15.770 3.285 16.110 3.620 ;
        RECT 18.010 3.285 18.350 3.620 ;
        RECT 20.250 3.285 20.590 3.620 ;
        RECT 22.545 2.640 22.775 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 23.950 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 23.950 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.015 ;
        RECT 2.430 0.300 2.770 0.635 ;
        RECT 4.670 0.300 5.010 0.635 ;
        RECT 6.910 0.300 7.250 0.635 ;
        RECT 9.150 0.300 9.490 0.635 ;
        RECT 11.390 0.300 11.730 0.635 ;
        RECT 13.630 0.300 13.970 0.635 ;
        RECT 15.870 0.300 16.210 0.635 ;
        RECT 18.110 0.300 18.450 0.635 ;
        RECT 20.350 0.300 20.690 0.635 ;
        RECT 22.645 0.300 22.875 1.015 ;
        RECT 0.000 -0.300 23.520 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__inv_20
MACRO gf180mcu_fd_sc_mcu7t5v0__invz_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__invz_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.052000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.410 1.700 2.425 2.120 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.526000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.740 1.560 9.400 2.375 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.072725 ;
    PORT
      LAYER Metal1 ;
        RECT 4.530 0.990 4.920 2.930 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 9.520 4.220 ;
        RECT 1.265 2.865 1.495 3.620 ;
        RECT 5.615 3.000 5.845 3.620 ;
        RECT 7.770 3.115 8.000 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 9.950 4.350 ;
        RECT -0.430 1.760 3.390 1.885 ;
        RECT 5.255 1.760 9.950 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 3.390 1.760 5.255 1.885 ;
        RECT -0.430 -0.430 9.950 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.760 ;
        RECT 5.930 0.300 6.160 0.905 ;
        RECT 7.770 0.300 8.000 0.815 ;
        RECT 0.000 -0.300 9.520 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.635 0.475 3.390 ;
        RECT 2.285 3.160 5.385 3.390 ;
        RECT 2.285 2.865 2.515 3.160 ;
        RECT 0.245 2.405 3.010 2.635 ;
        RECT 2.710 1.225 3.010 2.405 ;
        RECT 0.180 0.995 3.010 1.225 ;
        RECT 3.240 2.610 3.820 2.910 ;
        RECT 0.180 0.530 0.540 0.995 ;
        RECT 3.240 0.760 3.470 2.610 ;
        RECT 4.050 2.380 4.280 3.160 ;
        RECT 3.770 2.150 4.280 2.380 ;
        RECT 5.150 2.770 5.385 3.160 ;
        RECT 6.750 2.770 6.980 3.375 ;
        RECT 8.945 2.885 9.175 3.375 ;
        RECT 5.150 2.535 6.980 2.770 ;
        RECT 7.260 2.650 9.175 2.885 ;
        RECT 3.770 0.990 4.110 2.150 ;
        RECT 5.150 1.900 5.380 2.535 ;
        RECT 5.345 1.365 5.575 1.620 ;
        RECT 5.345 1.135 6.935 1.365 ;
        RECT 5.345 0.760 5.575 1.135 ;
        RECT 2.400 0.530 5.575 0.760 ;
        RECT 6.585 0.530 6.935 1.135 ;
        RECT 7.260 1.275 7.490 2.650 ;
        RECT 7.260 1.045 8.460 1.275 ;
        RECT 8.230 0.760 8.460 1.045 ;
        RECT 8.230 0.530 9.340 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__invz_1
MACRO gf180mcu_fd_sc_mcu7t5v0__invz_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__invz_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.410 1.625 1.590 2.125 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.082000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.405 1.640 8.775 2.190 ;
        RECT 7.405 1.160 7.770 1.640 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.040000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.880 1.660 7.175 2.800 ;
        RECT 6.795 0.530 7.175 1.660 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 9.520 4.220 ;
        RECT 1.465 2.815 1.805 3.620 ;
        RECT 5.925 2.890 6.155 3.620 ;
        RECT 7.965 2.980 8.195 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 9.950 4.350 ;
        RECT -0.430 1.760 3.400 1.885 ;
        RECT 4.520 1.760 9.950 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 3.400 1.760 4.520 1.885 ;
        RECT -0.430 -0.430 9.950 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.375 0.300 1.605 0.760 ;
        RECT 5.620 0.300 5.960 0.635 ;
        RECT 7.915 0.300 8.145 0.920 ;
        RECT 0.000 -0.300 9.520 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.500 2.585 0.730 3.380 ;
        RECT 2.445 3.125 5.135 3.355 ;
        RECT 0.500 2.355 3.210 2.585 ;
        RECT 1.840 2.035 3.210 2.355 ;
        RECT 1.840 1.225 2.070 2.035 ;
        RECT 3.555 1.805 3.790 2.890 ;
        RECT 0.255 0.990 2.070 1.225 ;
        RECT 2.985 1.575 3.790 1.805 ;
        RECT 0.255 0.570 0.485 0.990 ;
        RECT 2.985 0.885 3.215 1.575 ;
        RECT 4.020 1.555 4.250 3.125 ;
        RECT 4.905 2.465 5.135 3.125 ;
        RECT 6.385 3.070 7.735 3.300 ;
        RECT 6.385 2.660 6.615 3.070 ;
        RECT 5.415 2.425 6.615 2.660 ;
        RECT 7.505 2.750 7.735 3.070 ;
        RECT 9.020 2.750 9.285 3.380 ;
        RECT 7.505 2.520 9.285 2.750 ;
        RECT 5.415 1.915 5.645 2.425 ;
        RECT 5.875 1.965 6.650 2.195 ;
        RECT 5.875 1.555 6.105 1.965 ;
        RECT 4.020 1.345 6.105 1.555 ;
        RECT 3.770 1.325 6.105 1.345 ;
        RECT 3.770 0.990 4.250 1.325 ;
        RECT 6.335 1.095 6.565 1.640 ;
        RECT 2.495 0.760 3.215 0.885 ;
        RECT 5.160 0.865 6.565 1.095 ;
        RECT 5.160 0.760 5.390 0.865 ;
        RECT 2.495 0.530 5.390 0.760 ;
        RECT 9.020 0.580 9.285 2.520 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__invz_2
MACRO gf180mcu_fd_sc_mcu7t5v0__invz_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__invz_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.880 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.660 1.650 1.600 2.150 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.039500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.530 1.790 6.110 2.125 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.920000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.410 2.660 9.750 3.165 ;
        RECT 11.450 2.750 11.790 3.165 ;
        RECT 11.450 2.660 12.760 2.750 ;
        RECT 9.410 2.425 12.760 2.660 ;
        RECT 12.265 1.100 12.760 2.425 ;
        RECT 10.025 0.865 12.760 1.100 ;
        RECT 10.025 0.615 10.255 0.865 ;
        RECT 12.265 0.610 12.760 0.865 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 12.880 4.220 ;
        RECT 1.565 3.065 1.795 3.620 ;
        RECT 6.085 3.285 6.425 3.620 ;
        RECT 8.335 2.760 8.565 3.620 ;
        RECT 10.485 3.165 10.715 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 13.310 4.350 ;
        RECT -0.430 1.760 3.445 1.885 ;
        RECT 5.420 1.760 13.310 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 3.445 1.760 5.420 1.885 ;
        RECT -0.430 -0.430 13.310 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.420 0.300 1.650 0.760 ;
        RECT 6.130 0.300 6.470 0.635 ;
        RECT 8.725 0.300 8.955 0.900 ;
        RECT 11.090 0.300 11.430 0.635 ;
        RECT 0.000 -0.300 12.880 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.545 2.790 0.775 3.305 ;
        RECT 2.530 3.155 5.715 3.390 ;
        RECT 0.545 2.495 3.255 2.790 ;
        RECT 1.860 2.035 3.255 2.495 ;
        RECT 1.860 1.225 2.090 2.035 ;
        RECT 3.600 1.805 3.835 2.890 ;
        RECT 0.300 0.990 2.090 1.225 ;
        RECT 3.030 1.575 3.835 1.805 ;
        RECT 0.300 0.675 0.530 0.990 ;
        RECT 3.030 0.885 3.260 1.575 ;
        RECT 4.065 1.345 4.295 3.155 ;
        RECT 5.485 3.055 5.715 3.155 ;
        RECT 5.025 2.590 5.255 2.870 ;
        RECT 5.485 2.825 8.105 3.055 ;
        RECT 5.025 2.355 6.975 2.590 ;
        RECT 6.745 1.560 6.975 2.355 ;
        RECT 7.875 2.195 8.105 2.825 ;
        RECT 7.875 1.960 11.365 2.195 ;
        RECT 3.815 0.990 4.295 1.345 ;
        RECT 5.120 1.555 6.975 1.560 ;
        RECT 5.120 1.325 7.970 1.555 ;
        RECT 8.200 1.365 11.870 1.595 ;
        RECT 5.120 1.220 5.350 1.325 ;
        RECT 4.700 0.990 5.350 1.220 ;
        RECT 8.200 1.095 8.430 1.365 ;
        RECT 2.540 0.760 3.260 0.885 ;
        RECT 5.580 0.865 8.430 1.095 ;
        RECT 5.580 0.760 5.810 0.865 ;
        RECT 2.540 0.530 5.810 0.760 ;
        RECT 7.395 0.530 7.625 0.865 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__invz_3
MACRO gf180mcu_fd_sc_mcu7t5v0__invz_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__invz_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.440 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.370 1.760 1.620 2.150 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.039500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.475 1.790 6.070 2.135 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.080000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.110 2.660 9.410 3.380 ;
        RECT 11.190 2.660 11.420 3.380 ;
        RECT 9.110 2.425 11.420 2.660 ;
        RECT 10.730 1.100 11.110 2.425 ;
        RECT 9.400 0.865 11.870 1.100 ;
        RECT 9.400 0.715 9.630 0.865 ;
        RECT 11.640 0.710 11.870 0.865 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 13.440 4.220 ;
        RECT 1.455 3.285 1.795 3.620 ;
        RECT 5.985 3.285 6.325 3.620 ;
        RECT 8.075 2.815 8.415 3.620 ;
        RECT 10.170 3.020 10.400 3.620 ;
        RECT 12.210 2.565 12.440 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 13.870 4.350 ;
        RECT -0.430 1.760 3.390 1.885 ;
        RECT 5.235 1.760 13.870 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 3.390 1.760 5.235 1.885 ;
        RECT -0.430 -0.430 13.870 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 0.760 ;
        RECT 5.985 0.300 6.325 0.635 ;
        RECT 8.225 0.300 8.565 0.635 ;
        RECT 10.465 0.300 10.805 0.635 ;
        RECT 12.760 0.300 12.990 1.060 ;
        RECT 0.000 -0.300 13.440 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.490 2.740 0.720 3.380 ;
        RECT 2.475 3.125 5.625 3.355 ;
        RECT 4.010 3.120 5.625 3.125 ;
        RECT 0.490 2.510 2.100 2.740 ;
        RECT 1.870 2.320 2.100 2.510 ;
        RECT 1.870 2.085 3.260 2.320 ;
        RECT 1.870 1.225 2.100 2.085 ;
        RECT 3.545 1.805 3.780 2.890 ;
        RECT 0.245 0.990 2.100 1.225 ;
        RECT 2.975 1.575 3.780 1.805 ;
        RECT 0.245 0.670 0.475 0.990 ;
        RECT 2.975 0.885 3.205 1.575 ;
        RECT 4.010 1.345 4.240 3.120 ;
        RECT 5.395 3.055 5.625 3.120 ;
        RECT 7.110 3.055 7.340 3.380 ;
        RECT 4.890 2.595 5.120 2.890 ;
        RECT 5.395 2.825 7.340 3.055 ;
        RECT 4.890 2.365 6.830 2.595 ;
        RECT 6.600 2.125 6.830 2.365 ;
        RECT 7.110 2.585 7.340 2.825 ;
        RECT 7.110 2.355 8.565 2.585 ;
        RECT 8.335 2.195 8.565 2.355 ;
        RECT 6.600 1.730 7.940 2.125 ;
        RECT 8.335 1.960 9.950 2.195 ;
        RECT 6.600 1.560 6.830 1.730 ;
        RECT 3.760 0.990 4.240 1.345 ;
        RECT 4.935 1.325 6.830 1.560 ;
        RECT 8.335 1.365 10.125 1.595 ;
        RECT 4.935 1.220 5.165 1.325 ;
        RECT 4.515 0.990 5.165 1.220 ;
        RECT 8.335 1.095 8.565 1.365 ;
        RECT 2.485 0.760 3.205 0.885 ;
        RECT 5.395 0.865 8.565 1.095 ;
        RECT 5.395 0.760 5.625 0.865 ;
        RECT 2.485 0.530 5.625 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__invz_4
MACRO gf180mcu_fd_sc_mcu7t5v0__invz_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__invz_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.840 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.370 1.770 1.625 2.150 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.073000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.570 1.785 7.720 2.150 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.267600 ;
    PORT
      LAYER Metal1 ;
        RECT 13.505 2.830 13.745 3.380 ;
        RECT 15.600 2.830 15.830 3.380 ;
        RECT 17.640 2.830 17.870 3.380 ;
        RECT 19.680 2.830 19.910 3.380 ;
        RECT 13.505 2.530 19.910 2.830 ;
        RECT 16.850 1.155 17.340 2.530 ;
        RECT 15.740 1.135 18.315 1.155 ;
        RECT 13.510 0.865 20.460 1.135 ;
        RECT 13.510 0.630 13.740 0.865 ;
        RECT 15.750 0.635 15.980 0.865 ;
        RECT 17.990 0.635 18.220 0.865 ;
        RECT 20.230 0.635 20.460 0.865 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 21.840 4.220 ;
        RECT 1.535 3.285 1.880 3.620 ;
        RECT 4.955 3.445 5.295 3.620 ;
        RECT 7.555 3.445 7.915 3.620 ;
        RECT 10.100 2.665 10.330 3.620 ;
        RECT 12.340 2.665 12.570 3.620 ;
        RECT 14.580 3.230 14.810 3.620 ;
        RECT 16.620 3.230 16.850 3.620 ;
        RECT 18.660 3.230 18.890 3.620 ;
        RECT 20.700 2.530 20.930 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 22.270 4.350 ;
        RECT -0.430 1.760 3.405 1.885 ;
        RECT 7.235 1.760 22.270 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 3.405 1.760 7.235 1.885 ;
        RECT -0.430 -0.430 22.270 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.380 0.300 1.610 0.760 ;
        RECT 5.010 0.300 5.295 0.530 ;
        RECT 7.855 0.300 8.195 0.635 ;
        RECT 10.150 0.300 10.380 0.865 ;
        RECT 12.390 0.300 12.620 0.865 ;
        RECT 14.575 0.300 14.915 0.635 ;
        RECT 16.815 0.300 17.155 0.635 ;
        RECT 19.055 0.300 19.395 0.635 ;
        RECT 21.350 0.300 21.580 1.015 ;
        RECT 0.000 -0.300 21.840 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.575 2.800 0.805 3.380 ;
        RECT 2.520 3.215 4.725 3.355 ;
        RECT 5.525 3.215 7.325 3.355 ;
        RECT 2.520 3.125 9.365 3.215 ;
        RECT 4.095 3.055 9.365 3.125 ;
        RECT 4.095 2.985 5.875 3.055 ;
        RECT 6.810 2.985 9.365 3.055 ;
        RECT 0.575 2.570 2.185 2.800 ;
        RECT 1.955 2.320 2.185 2.570 ;
        RECT 1.955 2.090 3.345 2.320 ;
        RECT 1.955 1.225 2.185 2.090 ;
        RECT 3.635 1.805 3.865 2.890 ;
        RECT 0.260 0.990 2.185 1.225 ;
        RECT 2.990 1.575 3.865 1.805 ;
        RECT 0.260 0.675 0.490 0.990 ;
        RECT 2.990 0.885 3.220 1.575 ;
        RECT 4.095 1.345 4.325 2.985 ;
        RECT 6.105 2.755 6.580 2.780 ;
        RECT 6.105 2.525 8.730 2.755 ;
        RECT 8.500 1.955 8.730 2.525 ;
        RECT 9.025 2.415 9.365 2.985 ;
        RECT 11.220 2.415 11.450 3.260 ;
        RECT 9.025 2.195 12.620 2.415 ;
        RECT 9.025 2.185 16.325 2.195 ;
        RECT 12.390 1.960 16.325 2.185 ;
        RECT 18.165 1.960 20.460 2.195 ;
        RECT 8.500 1.625 12.145 1.955 ;
        RECT 8.500 1.555 8.730 1.625 ;
        RECT 3.775 1.115 4.325 1.345 ;
        RECT 6.515 1.325 8.730 1.555 ;
        RECT 12.390 1.365 15.480 1.595 ;
        RECT 18.505 1.365 21.140 1.595 ;
        RECT 12.390 1.325 12.620 1.365 ;
        RECT 3.775 0.990 4.135 1.115 ;
        RECT 6.515 0.990 6.935 1.325 ;
        RECT 9.405 1.095 12.620 1.325 ;
        RECT 2.500 0.760 3.220 0.885 ;
        RECT 4.550 0.760 6.000 0.990 ;
        RECT 7.165 0.865 9.635 1.095 ;
        RECT 7.165 0.760 7.395 0.865 ;
        RECT 2.500 0.530 4.780 0.760 ;
        RECT 5.770 0.530 7.395 0.760 ;
        RECT 9.030 0.530 9.260 0.865 ;
        RECT 11.270 0.530 11.500 1.095 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__invz_8
MACRO gf180mcu_fd_sc_mcu7t5v0__invz_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__invz_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.240 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.370 1.770 1.590 2.150 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.118500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.615 1.770 8.475 2.150 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.594000 ;
    PORT
      LAYER Metal1 ;
        RECT 17.445 2.860 17.675 3.380 ;
        RECT 19.585 2.860 19.815 3.380 ;
        RECT 21.825 2.860 22.055 3.380 ;
        RECT 23.965 2.860 24.195 3.380 ;
        RECT 26.005 2.860 26.235 3.380 ;
        RECT 28.045 2.860 28.280 3.380 ;
        RECT 17.445 2.460 28.280 2.860 ;
        RECT 23.040 1.265 23.440 2.460 ;
        RECT 20.750 1.135 26.610 1.265 ;
        RECT 17.120 0.865 28.880 1.135 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 30.240 4.220 ;
        RECT 1.630 3.130 1.860 3.620 ;
        RECT 6.400 3.445 6.740 3.620 ;
        RECT 9.815 3.100 10.045 3.620 ;
        RECT 12.020 2.590 12.360 3.620 ;
        RECT 14.060 2.590 14.400 3.620 ;
        RECT 16.170 2.590 16.510 3.620 ;
        RECT 18.465 3.230 18.695 3.620 ;
        RECT 20.705 3.230 20.935 3.620 ;
        RECT 22.945 3.230 23.175 3.620 ;
        RECT 24.985 3.230 25.215 3.620 ;
        RECT 27.025 3.230 27.255 3.620 ;
        RECT 29.065 2.530 29.295 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 30.670 4.350 ;
        RECT -0.430 1.760 3.440 1.885 ;
        RECT 8.440 1.760 30.670 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 3.440 1.760 8.440 1.885 ;
        RECT -0.430 -0.430 30.670 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.415 0.300 1.645 0.760 ;
        RECT 6.150 0.300 6.510 0.475 ;
        RECT 9.270 0.300 9.630 0.475 ;
        RECT 11.795 0.300 12.025 0.930 ;
        RECT 14.035 0.300 14.265 0.930 ;
        RECT 16.275 0.300 16.505 0.930 ;
        RECT 18.460 0.300 18.800 0.635 ;
        RECT 20.700 0.300 21.040 0.635 ;
        RECT 22.940 0.300 23.280 0.635 ;
        RECT 25.180 0.300 25.520 0.635 ;
        RECT 27.225 0.300 27.760 0.635 ;
        RECT 29.715 0.300 29.945 0.915 ;
        RECT 0.000 -0.300 30.240 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.610 2.865 0.840 3.380 ;
        RECT 2.595 3.215 6.170 3.355 ;
        RECT 6.970 3.215 9.490 3.355 ;
        RECT 2.595 3.125 9.490 3.215 ;
        RECT 4.130 3.010 9.490 3.125 ;
        RECT 0.610 2.570 2.165 2.865 ;
        RECT 1.935 2.320 2.165 2.570 ;
        RECT 1.935 2.090 3.375 2.320 ;
        RECT 1.935 1.225 2.165 2.090 ;
        RECT 3.670 1.860 3.900 2.890 ;
        RECT 0.295 0.990 2.165 1.225 ;
        RECT 3.025 1.630 3.900 1.860 ;
        RECT 0.295 0.715 0.525 0.990 ;
        RECT 3.025 0.885 3.255 1.630 ;
        RECT 4.130 1.400 4.360 3.010 ;
        RECT 5.940 2.985 7.200 3.010 ;
        RECT 9.260 2.840 9.490 3.010 ;
        RECT 11.055 2.840 11.285 3.380 ;
        RECT 5.150 2.755 5.665 2.780 ;
        RECT 7.430 2.755 9.000 2.780 ;
        RECT 5.150 2.525 9.000 2.755 ;
        RECT 9.260 2.610 11.285 2.840 ;
        RECT 3.810 0.990 4.360 1.400 ;
        RECT 8.770 1.900 9.000 2.525 ;
        RECT 11.055 2.360 11.285 2.610 ;
        RECT 13.095 2.360 13.325 3.380 ;
        RECT 15.135 2.360 15.365 3.380 ;
        RECT 11.055 2.195 16.505 2.360 ;
        RECT 11.055 2.130 22.650 2.195 ;
        RECT 16.275 1.960 22.650 2.130 ;
        RECT 24.405 1.960 28.840 2.195 ;
        RECT 8.770 1.650 15.965 1.900 ;
        RECT 8.770 1.395 9.000 1.650 ;
        RECT 16.275 1.420 20.475 1.595 ;
        RECT 4.590 1.165 9.000 1.395 ;
        RECT 11.055 1.365 20.475 1.420 ;
        RECT 26.860 1.365 29.485 1.595 ;
        RECT 11.055 1.190 16.505 1.365 ;
        RECT 4.590 0.990 4.950 1.165 ;
        RECT 7.710 0.990 8.070 1.165 ;
        RECT 11.055 0.935 11.285 1.190 ;
        RECT 2.535 0.760 3.255 0.885 ;
        RECT 5.690 0.760 7.155 0.935 ;
        RECT 8.555 0.760 11.285 0.935 ;
        RECT 2.535 0.705 11.285 0.760 ;
        RECT 2.535 0.530 5.920 0.705 ;
        RECT 6.925 0.530 8.785 0.705 ;
        RECT 12.915 0.580 13.145 1.190 ;
        RECT 15.155 0.580 15.385 1.190 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__invz_12
MACRO gf180mcu_fd_sc_mcu7t5v0__invz_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__invz_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 39.200 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.370 1.770 1.590 2.150 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.130 1.770 9.850 2.150 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.205000 ;
    PORT
      LAYER Metal1 ;
        RECT 21.820 3.005 22.050 3.380 ;
        RECT 24.025 3.005 24.255 3.380 ;
        RECT 26.255 3.005 26.485 3.380 ;
        RECT 28.510 3.005 28.740 3.380 ;
        RECT 30.755 3.005 30.985 3.380 ;
        RECT 32.975 3.005 33.205 3.380 ;
        RECT 35.225 3.005 35.455 3.380 ;
        RECT 37.500 3.005 37.785 3.380 ;
        RECT 21.820 2.425 37.785 3.005 ;
        RECT 28.950 1.445 29.850 2.425 ;
        RECT 25.240 1.135 34.285 1.445 ;
        RECT 21.755 0.865 37.785 1.135 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 39.200 4.220 ;
        RECT 1.630 3.285 1.970 3.620 ;
        RECT 5.045 3.445 5.385 3.620 ;
        RECT 8.155 3.445 8.515 3.620 ;
        RECT 11.350 2.700 11.580 3.620 ;
        RECT 13.760 2.700 13.990 3.620 ;
        RECT 15.995 2.700 16.225 3.620 ;
        RECT 18.330 2.700 18.560 3.620 ;
        RECT 20.680 2.700 20.910 3.620 ;
        RECT 22.835 3.285 23.175 3.620 ;
        RECT 25.080 3.285 25.420 3.620 ;
        RECT 27.330 3.285 27.670 3.620 ;
        RECT 29.570 3.285 29.910 3.620 ;
        RECT 31.810 3.285 32.150 3.620 ;
        RECT 34.050 3.285 34.390 3.620 ;
        RECT 36.285 3.285 36.625 3.620 ;
        RECT 38.520 2.530 38.750 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 39.630 4.350 ;
        RECT -0.430 1.760 3.495 1.885 ;
        RECT 10.445 1.760 39.630 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 3.495 1.760 10.445 1.885 ;
        RECT -0.430 -0.430 39.630 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.470 0.300 1.700 0.760 ;
        RECT 5.100 0.300 5.385 0.530 ;
        RECT 8.155 0.300 8.515 0.475 ;
        RECT 11.275 0.300 11.635 0.475 ;
        RECT 13.800 0.300 14.030 0.870 ;
        RECT 16.040 0.300 16.270 0.870 ;
        RECT 18.280 0.300 18.510 0.870 ;
        RECT 20.700 0.300 20.930 0.870 ;
        RECT 22.885 0.300 23.225 0.635 ;
        RECT 25.125 0.300 25.465 0.635 ;
        RECT 27.365 0.300 27.705 0.635 ;
        RECT 29.605 0.300 29.945 0.635 ;
        RECT 31.845 0.300 32.185 0.635 ;
        RECT 34.085 0.300 34.425 0.635 ;
        RECT 36.325 0.300 36.665 0.635 ;
        RECT 38.620 0.300 38.850 1.015 ;
        RECT 0.000 -0.300 39.200 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.665 2.800 0.895 3.380 ;
        RECT 2.590 3.215 4.815 3.350 ;
        RECT 5.615 3.215 7.615 3.355 ;
        RECT 8.855 3.215 11.045 3.355 ;
        RECT 2.590 3.120 11.045 3.215 ;
        RECT 4.185 3.010 11.045 3.120 ;
        RECT 4.185 2.985 5.845 3.010 ;
        RECT 7.385 2.985 9.085 3.010 ;
        RECT 0.665 2.570 3.375 2.800 ;
        RECT 2.045 2.035 3.375 2.570 ;
        RECT 2.045 1.225 2.275 2.035 ;
        RECT 3.725 1.805 3.955 2.890 ;
        RECT 0.350 0.990 2.275 1.225 ;
        RECT 3.080 1.575 3.955 1.805 ;
        RECT 0.350 0.675 0.580 0.990 ;
        RECT 3.080 0.885 3.310 1.575 ;
        RECT 4.185 1.345 4.415 2.985 ;
        RECT 6.310 2.755 7.125 2.780 ;
        RECT 9.315 2.755 10.405 2.780 ;
        RECT 6.310 2.525 10.405 2.755 ;
        RECT 10.175 1.960 10.405 2.525 ;
        RECT 10.815 2.425 11.045 3.010 ;
        RECT 12.630 2.425 12.860 3.380 ;
        RECT 14.880 2.425 15.110 3.380 ;
        RECT 17.125 2.425 17.355 3.380 ;
        RECT 19.520 2.425 19.750 3.380 ;
        RECT 10.815 2.195 20.930 2.425 ;
        RECT 10.815 2.190 28.145 2.195 ;
        RECT 20.700 1.960 28.145 2.190 ;
        RECT 32.315 1.960 38.300 2.195 ;
        RECT 10.175 1.630 20.325 1.960 ;
        RECT 10.175 1.420 10.415 1.630 ;
        RECT 3.865 1.115 4.415 1.345 ;
        RECT 6.595 1.190 10.415 1.420 ;
        RECT 20.700 1.365 24.785 1.595 ;
        RECT 34.765 1.365 38.300 1.595 ;
        RECT 20.700 1.330 20.930 1.365 ;
        RECT 3.865 0.990 4.225 1.115 ;
        RECT 6.595 0.990 6.955 1.190 ;
        RECT 9.715 0.990 10.415 1.190 ;
        RECT 13.025 1.100 20.930 1.330 ;
        RECT 2.590 0.760 3.310 0.885 ;
        RECT 4.640 0.760 6.365 0.990 ;
        RECT 13.025 0.960 13.255 1.100 ;
        RECT 7.185 0.760 9.485 0.960 ;
        RECT 10.815 0.760 13.255 0.960 ;
        RECT 2.590 0.530 4.870 0.760 ;
        RECT 6.135 0.730 13.255 0.760 ;
        RECT 6.135 0.530 7.415 0.730 ;
        RECT 9.255 0.530 11.045 0.730 ;
        RECT 14.920 0.530 15.150 1.100 ;
        RECT 17.160 0.530 17.390 1.100 ;
        RECT 19.580 0.530 19.810 1.100 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__invz_16
MACRO gf180mcu_fd_sc_mcu7t5v0__latq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.200 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 1.240 4.430 1.560 ;
        RECT 4.000 0.550 4.430 1.240 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.736000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.770 2.120 2.150 2.750 ;
        RECT 0.825 1.800 2.150 2.120 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 9.605 0.530 9.960 3.380 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 11.200 4.220 ;
        RECT 1.265 2.660 1.495 3.620 ;
        RECT 3.485 3.085 3.715 3.620 ;
        RECT 7.765 2.655 7.995 3.620 ;
        RECT 10.625 2.530 10.855 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 11.630 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 11.630 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 0.815 ;
        RECT 3.385 0.300 3.615 0.825 ;
        RECT 7.765 0.300 7.995 0.895 ;
        RECT 10.725 0.300 10.955 1.160 ;
        RECT 0.000 -0.300 11.200 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 1.390 0.530 3.390 ;
        RECT 2.610 2.085 2.895 3.390 ;
        RECT 5.100 3.140 6.505 3.370 ;
        RECT 3.125 2.335 5.100 2.565 ;
        RECT 5.755 2.085 5.985 2.810 ;
        RECT 2.610 1.855 5.985 2.085 ;
        RECT 0.190 1.160 2.360 1.390 ;
        RECT 0.190 0.530 0.530 1.160 ;
        RECT 2.610 0.530 2.950 1.855 ;
        RECT 4.785 1.010 5.015 1.855 ;
        RECT 6.275 1.475 6.505 3.140 ;
        RECT 8.785 2.305 9.035 3.225 ;
        RECT 7.025 2.075 9.170 2.305 ;
        RECT 6.275 1.245 8.580 1.475 ;
        RECT 6.275 0.760 6.505 1.245 ;
        RECT 5.200 0.530 6.505 0.760 ;
        RECT 8.830 0.530 9.170 2.075 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latq_1
MACRO gf180mcu_fd_sc_mcu7t5v0__latq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.320 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 1.240 4.430 1.560 ;
        RECT 4.000 0.550 4.430 1.240 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.736000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.770 2.120 2.150 2.750 ;
        RECT 0.825 1.800 2.150 2.120 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.060800 ;
    PORT
      LAYER Metal1 ;
        RECT 10.660 0.530 11.080 3.380 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 12.320 4.220 ;
        RECT 1.365 3.050 1.595 3.620 ;
        RECT 3.485 3.085 3.715 3.620 ;
        RECT 7.410 2.805 7.750 3.620 ;
        RECT 9.705 2.530 9.935 3.620 ;
        RECT 11.745 2.530 11.975 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 12.750 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.750 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 0.815 ;
        RECT 3.385 0.300 3.615 0.825 ;
        RECT 7.765 0.300 7.995 0.895 ;
        RECT 9.605 0.300 9.835 1.055 ;
        RECT 11.845 0.300 12.075 1.055 ;
        RECT 0.000 -0.300 12.320 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 1.390 0.575 3.390 ;
        RECT 2.610 2.085 2.895 3.390 ;
        RECT 5.100 3.140 6.505 3.370 ;
        RECT 3.125 2.335 5.100 2.565 ;
        RECT 5.755 2.085 5.985 2.810 ;
        RECT 2.610 1.855 5.985 2.085 ;
        RECT 0.190 1.160 2.360 1.390 ;
        RECT 0.190 0.530 0.575 1.160 ;
        RECT 2.610 0.530 2.950 1.855 ;
        RECT 4.785 1.010 5.015 1.855 ;
        RECT 6.275 1.475 6.505 3.140 ;
        RECT 8.485 2.305 8.715 3.225 ;
        RECT 6.820 2.075 9.170 2.305 ;
        RECT 6.275 1.245 8.580 1.475 ;
        RECT 6.275 0.760 6.505 1.245 ;
        RECT 5.200 0.530 6.505 0.760 ;
        RECT 8.830 0.530 9.170 2.075 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latq_2
MACRO gf180mcu_fd_sc_mcu7t5v0__latq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.680 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 1.240 4.430 1.560 ;
        RECT 4.000 0.550 4.430 1.240 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.736000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 2.120 2.150 2.750 ;
        RECT 0.825 1.800 2.150 2.120 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.121600 ;
    PORT
      LAYER Metal1 ;
        RECT 11.240 2.120 11.700 3.380 ;
        RECT 13.280 2.120 13.880 3.380 ;
        RECT 11.240 1.800 13.880 2.120 ;
        RECT 11.240 0.530 11.700 1.800 ;
        RECT 13.280 0.530 13.880 1.800 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 15.680 4.220 ;
        RECT 1.365 3.050 1.595 3.620 ;
        RECT 3.485 3.085 3.715 3.620 ;
        RECT 7.705 2.805 8.050 3.620 ;
        RECT 10.225 2.530 10.455 3.620 ;
        RECT 12.265 2.530 12.495 3.620 ;
        RECT 14.305 2.530 14.535 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 16.110 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 16.110 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 0.815 ;
        RECT 3.385 0.300 3.615 0.825 ;
        RECT 7.765 0.300 7.995 0.895 ;
        RECT 10.225 0.300 10.455 1.055 ;
        RECT 12.465 0.300 12.695 1.055 ;
        RECT 14.705 0.300 14.935 1.055 ;
        RECT 0.000 -0.300 15.680 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 1.390 0.575 3.390 ;
        RECT 2.610 2.085 2.895 3.390 ;
        RECT 5.100 3.140 6.505 3.370 ;
        RECT 3.125 2.335 5.100 2.565 ;
        RECT 5.755 2.085 5.985 2.810 ;
        RECT 2.610 1.855 5.985 2.085 ;
        RECT 0.190 1.160 2.360 1.390 ;
        RECT 0.190 0.530 0.575 1.160 ;
        RECT 2.610 0.530 2.950 1.855 ;
        RECT 4.785 1.010 5.015 1.855 ;
        RECT 6.275 1.475 6.505 3.140 ;
        RECT 8.785 2.305 9.015 3.225 ;
        RECT 7.120 2.075 9.170 2.305 ;
        RECT 6.275 1.245 8.580 1.475 ;
        RECT 6.275 0.760 6.505 1.245 ;
        RECT 5.200 0.530 6.505 0.760 ;
        RECT 8.830 0.530 9.170 2.075 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latq_4
MACRO gf180mcu_fd_sc_mcu7t5v0__latrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latrnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.320 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.285 1.240 3.310 1.630 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.293500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.760 1.045 2.055 1.275 ;
        RECT 5.160 1.265 5.475 2.135 ;
        RECT 1.825 1.000 2.055 1.045 ;
        RECT 3.675 1.035 5.475 1.265 ;
        RECT 3.675 1.000 3.905 1.035 ;
        RECT 1.825 0.680 3.905 1.000 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.789000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 2.595 5.935 2.680 ;
        RECT 2.380 2.365 5.935 2.595 ;
        RECT 5.705 1.795 5.935 2.365 ;
        RECT 5.705 1.565 7.000 1.795 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 11.530 2.530 12.190 3.380 ;
        RECT 11.880 1.120 12.190 2.530 ;
        RECT 11.310 0.600 12.190 1.120 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 12.320 4.220 ;
        RECT 1.265 2.655 1.495 3.620 ;
        RECT 2.970 3.285 3.310 3.620 ;
        RECT 6.960 3.285 7.300 3.620 ;
        RECT 10.510 2.815 10.850 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 12.750 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.750 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 0.815 ;
        RECT 7.325 0.300 7.555 0.875 ;
        RECT 10.285 0.300 10.515 1.075 ;
        RECT 0.000 -0.300 12.320 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 2.135 0.475 3.310 ;
        RECT 2.005 3.055 2.235 3.390 ;
        RECT 3.560 3.105 6.445 3.335 ;
        RECT 3.560 3.055 3.790 3.105 ;
        RECT 2.005 2.825 3.790 3.055 ;
        RECT 6.195 3.055 6.445 3.105 ;
        RECT 6.195 2.825 8.115 3.055 ;
        RECT 6.165 2.195 7.545 2.535 ;
        RECT 7.775 2.250 8.115 2.825 ;
        RECT 0.190 1.905 4.640 2.135 ;
        RECT 7.315 2.020 7.545 2.195 ;
        RECT 8.345 2.020 8.575 3.390 ;
        RECT 9.165 2.570 9.395 3.250 ;
        RECT 9.165 2.340 10.575 2.570 ;
        RECT 10.345 2.020 10.575 2.340 ;
        RECT 0.190 0.530 0.530 1.905 ;
        RECT 7.315 1.790 10.005 2.020 ;
        RECT 10.345 1.790 11.310 2.020 ;
        RECT 6.865 1.105 8.170 1.335 ;
        RECT 6.865 0.760 7.095 1.105 ;
        RECT 4.290 0.530 7.095 0.760 ;
        RECT 8.445 0.550 8.675 1.790 ;
        RECT 10.345 1.535 10.575 1.790 ;
        RECT 9.165 1.305 10.575 1.535 ;
        RECT 9.165 0.735 9.395 1.305 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latrnq_1
MACRO gf180mcu_fd_sc_mcu7t5v0__latrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latrnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.440 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.285 1.240 3.310 1.630 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.293500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.760 1.045 2.055 1.275 ;
        RECT 5.160 1.265 5.475 2.135 ;
        RECT 1.825 1.000 2.055 1.045 ;
        RECT 3.675 1.035 5.475 1.265 ;
        RECT 3.675 1.000 3.905 1.035 ;
        RECT 1.825 0.680 3.905 1.000 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.789000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 2.595 5.935 2.680 ;
        RECT 2.380 2.365 5.935 2.595 ;
        RECT 5.705 1.795 5.935 2.365 ;
        RECT 5.705 1.565 7.000 1.795 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.060800 ;
    PORT
      LAYER Metal1 ;
        RECT 11.530 2.530 12.220 3.380 ;
        RECT 11.900 1.120 12.220 2.530 ;
        RECT 11.310 0.600 12.220 1.120 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 13.440 4.220 ;
        RECT 1.265 2.655 1.495 3.620 ;
        RECT 2.970 3.285 3.310 3.620 ;
        RECT 6.960 3.285 7.300 3.620 ;
        RECT 10.510 2.815 10.850 3.620 ;
        RECT 12.605 2.530 12.835 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 13.870 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.870 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 0.815 ;
        RECT 7.325 0.300 7.555 0.875 ;
        RECT 10.285 0.300 10.515 1.075 ;
        RECT 12.705 0.300 12.935 1.075 ;
        RECT 0.000 -0.300 13.440 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 2.135 0.475 3.310 ;
        RECT 2.005 3.055 2.235 3.390 ;
        RECT 3.560 3.105 6.445 3.335 ;
        RECT 3.560 3.055 3.790 3.105 ;
        RECT 2.005 2.825 3.790 3.055 ;
        RECT 6.195 3.055 6.445 3.105 ;
        RECT 6.195 2.825 8.115 3.055 ;
        RECT 6.165 2.195 7.545 2.535 ;
        RECT 7.775 2.250 8.115 2.825 ;
        RECT 0.190 1.905 4.640 2.135 ;
        RECT 7.315 2.020 7.545 2.195 ;
        RECT 8.345 2.020 8.575 3.390 ;
        RECT 9.165 2.570 9.395 3.250 ;
        RECT 9.165 2.340 10.575 2.570 ;
        RECT 10.345 2.030 10.575 2.340 ;
        RECT 0.190 0.530 0.530 1.905 ;
        RECT 7.315 1.790 9.890 2.020 ;
        RECT 6.865 1.105 8.170 1.335 ;
        RECT 6.865 0.760 7.095 1.105 ;
        RECT 4.290 0.530 7.095 0.760 ;
        RECT 8.445 0.550 8.675 1.790 ;
        RECT 10.345 1.690 11.650 2.030 ;
        RECT 10.345 1.545 10.575 1.690 ;
        RECT 9.165 1.315 10.575 1.545 ;
        RECT 9.165 0.735 9.395 1.315 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latrnq_2
MACRO gf180mcu_fd_sc_mcu7t5v0__latrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latrnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.360 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.285 1.240 3.310 1.630 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.293500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.760 1.045 2.055 1.275 ;
        RECT 5.160 1.265 5.475 2.135 ;
        RECT 1.825 1.000 2.055 1.045 ;
        RECT 3.675 1.035 5.475 1.265 ;
        RECT 3.675 1.000 3.905 1.035 ;
        RECT 1.825 0.680 3.905 1.000 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.789000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 2.595 5.935 2.680 ;
        RECT 2.380 2.365 5.935 2.595 ;
        RECT 5.705 1.795 5.935 2.365 ;
        RECT 5.705 1.565 7.000 1.795 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.121600 ;
    PORT
      LAYER Metal1 ;
        RECT 13.205 2.585 13.435 3.380 ;
        RECT 15.240 2.585 15.590 3.380 ;
        RECT 13.205 2.355 15.590 2.585 ;
        RECT 15.240 1.560 15.590 2.355 ;
        RECT 13.105 1.240 15.590 1.560 ;
        RECT 13.105 0.550 13.335 1.240 ;
        RECT 15.240 0.550 15.590 1.240 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 17.360 4.220 ;
        RECT 1.265 2.655 1.495 3.620 ;
        RECT 2.970 3.285 3.310 3.620 ;
        RECT 6.960 3.285 7.300 3.620 ;
        RECT 9.565 2.655 9.795 3.620 ;
        RECT 11.650 2.815 11.990 3.620 ;
        RECT 14.170 2.815 14.510 3.620 ;
        RECT 16.210 2.625 16.550 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 17.790 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 17.790 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 0.815 ;
        RECT 7.325 0.300 7.555 0.875 ;
        RECT 9.565 0.300 9.795 0.890 ;
        RECT 11.805 0.300 12.035 0.890 ;
        RECT 14.225 0.300 14.455 0.890 ;
        RECT 16.465 0.300 16.695 0.930 ;
        RECT 0.000 -0.300 17.360 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 2.135 0.475 3.310 ;
        RECT 2.005 3.055 2.235 3.390 ;
        RECT 3.560 3.105 6.445 3.335 ;
        RECT 3.560 3.055 3.790 3.105 ;
        RECT 2.005 2.825 3.790 3.055 ;
        RECT 6.195 3.055 6.445 3.105 ;
        RECT 6.195 2.825 8.215 3.055 ;
        RECT 6.165 2.195 7.545 2.535 ;
        RECT 7.875 2.250 8.215 2.825 ;
        RECT 0.190 1.905 4.640 2.135 ;
        RECT 7.315 2.020 7.545 2.195 ;
        RECT 8.445 2.020 8.675 3.250 ;
        RECT 10.685 2.545 10.915 3.290 ;
        RECT 10.685 2.315 12.035 2.545 ;
        RECT 11.805 2.035 12.035 2.315 ;
        RECT 0.190 0.530 0.530 1.905 ;
        RECT 7.315 1.790 11.560 2.020 ;
        RECT 11.805 1.805 14.990 2.035 ;
        RECT 6.865 1.105 8.170 1.335 ;
        RECT 6.865 0.760 7.095 1.105 ;
        RECT 4.290 0.530 7.095 0.760 ;
        RECT 8.445 0.550 8.675 1.790 ;
        RECT 11.805 1.510 12.035 1.805 ;
        RECT 10.685 1.280 12.035 1.510 ;
        RECT 10.685 0.550 10.915 1.280 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latrnq_4
MACRO gf180mcu_fd_sc_mcu7t5v0__latrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latrsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.440 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.285 1.240 3.310 1.630 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.293500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.760 1.045 2.055 1.275 ;
        RECT 5.160 1.265 5.475 2.135 ;
        RECT 1.825 1.000 2.055 1.045 ;
        RECT 3.675 1.035 5.475 1.265 ;
        RECT 3.675 1.000 3.905 1.035 ;
        RECT 1.825 0.680 3.905 1.000 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.789000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 2.595 5.935 2.680 ;
        RECT 2.380 2.365 5.935 2.595 ;
        RECT 5.705 1.795 5.935 2.365 ;
        RECT 5.705 1.565 7.000 1.795 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.741500 ;
    PORT
      LAYER Metal1 ;
        RECT 9.010 1.085 9.400 2.355 ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 12.650 2.530 13.310 3.380 ;
        RECT 13.000 1.120 13.310 2.530 ;
        RECT 12.430 0.600 13.310 1.120 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 13.440 4.220 ;
        RECT 1.265 2.655 1.495 3.620 ;
        RECT 2.970 3.285 3.310 3.620 ;
        RECT 6.960 3.285 7.300 3.620 ;
        RECT 9.545 2.655 9.775 3.620 ;
        RECT 11.630 2.815 11.970 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 13.870 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.870 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 0.815 ;
        RECT 7.325 0.300 7.555 0.875 ;
        RECT 11.405 0.300 11.635 1.075 ;
        RECT 0.000 -0.300 13.440 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 2.135 0.475 3.310 ;
        RECT 2.005 3.055 2.235 3.390 ;
        RECT 3.560 3.105 6.445 3.335 ;
        RECT 3.560 3.055 3.790 3.105 ;
        RECT 2.005 2.825 3.790 3.055 ;
        RECT 6.195 3.055 6.445 3.105 ;
        RECT 6.195 2.825 8.115 3.055 ;
        RECT 6.165 2.195 7.545 2.535 ;
        RECT 7.775 2.250 8.115 2.825 ;
        RECT 0.190 1.905 4.640 2.135 ;
        RECT 7.315 2.020 7.545 2.195 ;
        RECT 8.525 2.020 8.755 3.390 ;
        RECT 10.285 2.570 10.515 3.250 ;
        RECT 10.285 2.340 11.695 2.570 ;
        RECT 11.465 2.020 11.695 2.340 ;
        RECT 0.190 0.530 0.530 1.905 ;
        RECT 7.315 1.790 8.755 2.020 ;
        RECT 6.865 1.105 8.115 1.335 ;
        RECT 6.865 0.760 7.095 1.105 ;
        RECT 4.290 0.530 7.095 0.760 ;
        RECT 8.525 0.835 8.755 1.790 ;
        RECT 9.760 1.790 11.125 2.020 ;
        RECT 11.465 1.790 12.430 2.020 ;
        RECT 9.760 0.835 9.990 1.790 ;
        RECT 11.465 1.535 11.695 1.790 ;
        RECT 8.525 0.605 9.990 0.835 ;
        RECT 10.285 1.305 11.695 1.535 ;
        RECT 10.285 0.735 10.515 1.305 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latrsnq_1
MACRO gf180mcu_fd_sc_mcu7t5v0__latrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latrsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.000 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.285 1.240 3.310 1.630 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.293500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.760 1.045 2.055 1.275 ;
        RECT 5.160 1.265 5.475 2.135 ;
        RECT 1.825 1.000 2.055 1.045 ;
        RECT 3.675 1.035 5.475 1.265 ;
        RECT 3.675 1.000 3.905 1.035 ;
        RECT 1.825 0.680 3.905 1.000 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.789000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 2.595 5.935 2.680 ;
        RECT 2.380 2.365 5.935 2.595 ;
        RECT 5.705 1.795 5.935 2.365 ;
        RECT 5.705 1.565 6.780 1.795 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.741500 ;
    PORT
      LAYER Metal1 ;
        RECT 8.840 1.085 9.400 2.355 ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.060800 ;
    PORT
      LAYER Metal1 ;
        RECT 12.380 2.380 12.760 3.380 ;
        RECT 12.380 2.150 13.340 2.380 ;
        RECT 12.980 1.365 13.340 2.150 ;
        RECT 12.380 1.135 13.340 1.365 ;
        RECT 12.380 0.545 12.760 1.135 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 14.000 4.220 ;
        RECT 1.265 2.655 1.495 3.620 ;
        RECT 2.970 3.285 3.310 3.620 ;
        RECT 6.960 3.285 7.300 3.620 ;
        RECT 9.345 2.655 9.575 3.620 ;
        RECT 11.210 2.630 11.550 3.620 ;
        RECT 13.350 2.630 13.690 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 14.430 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.430 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 0.815 ;
        RECT 7.325 0.300 7.555 0.875 ;
        RECT 11.265 0.300 11.495 0.885 ;
        RECT 13.505 0.300 13.735 0.885 ;
        RECT 0.000 -0.300 14.000 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 2.135 0.475 3.310 ;
        RECT 2.005 3.055 2.235 3.390 ;
        RECT 3.560 3.105 6.445 3.335 ;
        RECT 3.560 3.055 3.790 3.105 ;
        RECT 2.005 2.825 3.790 3.055 ;
        RECT 6.195 3.055 6.445 3.105 ;
        RECT 6.195 2.825 7.875 3.055 ;
        RECT 6.165 2.195 7.280 2.535 ;
        RECT 7.535 2.250 7.875 2.825 ;
        RECT 0.190 1.905 4.640 2.135 ;
        RECT 7.030 2.020 7.280 2.195 ;
        RECT 8.325 2.020 8.555 3.390 ;
        RECT 10.245 2.380 10.475 3.380 ;
        RECT 10.245 2.150 11.555 2.380 ;
        RECT 0.190 0.530 0.530 1.905 ;
        RECT 7.030 1.790 8.555 2.020 ;
        RECT 11.325 1.900 11.555 2.150 ;
        RECT 6.865 1.105 8.095 1.335 ;
        RECT 6.865 0.760 7.095 1.105 ;
        RECT 4.290 0.530 7.095 0.760 ;
        RECT 8.325 0.835 8.555 1.790 ;
        RECT 9.665 1.670 10.985 1.900 ;
        RECT 11.325 1.670 12.745 1.900 ;
        RECT 9.665 0.835 9.895 1.670 ;
        RECT 11.325 1.365 11.555 1.670 ;
        RECT 8.325 0.605 9.895 0.835 ;
        RECT 10.145 1.135 11.555 1.365 ;
        RECT 10.145 0.545 10.375 1.135 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latrsnq_2
MACRO gf180mcu_fd_sc_mcu7t5v0__latrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latrsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.360 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.285 1.240 3.310 1.630 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.293500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.760 1.045 2.055 1.275 ;
        RECT 5.160 1.265 5.475 2.135 ;
        RECT 1.825 1.000 2.055 1.045 ;
        RECT 3.675 1.035 5.475 1.265 ;
        RECT 3.675 1.000 3.905 1.035 ;
        RECT 1.825 0.680 3.905 1.000 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.789000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 2.595 5.935 2.680 ;
        RECT 2.380 2.365 5.935 2.595 ;
        RECT 5.705 1.795 5.935 2.365 ;
        RECT 5.705 1.565 6.780 1.795 ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.741500 ;
    PORT
      LAYER Metal1 ;
        RECT 8.840 1.085 9.400 2.355 ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.121600 ;
    PORT
      LAYER Metal1 ;
        RECT 13.540 2.570 13.900 3.380 ;
        RECT 15.645 2.570 16.140 3.380 ;
        RECT 13.540 2.340 16.680 2.570 ;
        RECT 16.350 1.465 16.680 2.340 ;
        RECT 13.505 1.160 16.680 1.465 ;
        RECT 13.505 0.545 13.735 1.160 ;
        RECT 15.745 0.545 15.975 1.160 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 17.360 4.220 ;
        RECT 1.265 2.655 1.495 3.620 ;
        RECT 2.970 3.285 3.310 3.620 ;
        RECT 6.960 3.285 7.300 3.620 ;
        RECT 9.345 2.655 9.575 3.620 ;
        RECT 10.245 2.530 10.475 3.620 ;
        RECT 12.380 2.815 12.720 3.620 ;
        RECT 14.570 2.815 14.910 3.620 ;
        RECT 16.610 2.815 16.950 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 17.790 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 17.790 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 0.815 ;
        RECT 7.325 0.300 7.555 0.875 ;
        RECT 10.145 0.300 10.375 0.885 ;
        RECT 12.385 0.300 12.615 0.885 ;
        RECT 14.625 0.300 14.855 0.885 ;
        RECT 16.865 0.300 17.095 0.885 ;
        RECT 0.000 -0.300 17.360 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 2.135 0.475 3.310 ;
        RECT 2.005 3.055 2.235 3.390 ;
        RECT 3.560 3.105 6.445 3.335 ;
        RECT 3.560 3.055 3.790 3.105 ;
        RECT 2.005 2.825 3.790 3.055 ;
        RECT 6.195 3.055 6.445 3.105 ;
        RECT 6.195 2.825 7.875 3.055 ;
        RECT 6.165 2.195 7.280 2.535 ;
        RECT 7.535 2.250 7.875 2.825 ;
        RECT 0.190 1.905 4.640 2.135 ;
        RECT 7.030 2.020 7.280 2.195 ;
        RECT 8.325 2.020 8.555 3.390 ;
        RECT 11.265 2.570 11.495 3.380 ;
        RECT 11.265 2.340 12.575 2.570 ;
        RECT 0.190 0.530 0.530 1.905 ;
        RECT 7.030 1.790 8.555 2.020 ;
        RECT 12.345 1.945 12.575 2.340 ;
        RECT 6.865 1.105 8.095 1.335 ;
        RECT 6.865 0.760 7.095 1.105 ;
        RECT 4.290 0.530 7.095 0.760 ;
        RECT 8.325 0.835 8.555 1.790 ;
        RECT 9.665 1.715 12.040 1.945 ;
        RECT 12.345 1.715 16.050 1.945 ;
        RECT 9.665 0.835 9.895 1.715 ;
        RECT 12.345 1.465 12.575 1.715 ;
        RECT 8.325 0.605 9.895 0.835 ;
        RECT 11.265 1.235 12.575 1.465 ;
        RECT 11.265 0.545 11.495 1.235 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latrsnq_4
MACRO gf180mcu_fd_sc_mcu7t5v0__latsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.760 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.965 1.790 3.270 2.120 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.293500 ;
    PORT
      LAYER Metal1 ;
        RECT 3.500 1.560 4.045 2.795 ;
        RECT 0.780 1.240 4.045 1.560 ;
    END
  END E
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.741500 ;
    PORT
      LAYER Metal1 ;
        RECT 5.040 1.800 7.380 2.120 ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 10.895 2.530 11.630 3.380 ;
        RECT 11.320 1.065 11.630 2.530 ;
        RECT 10.750 0.600 11.630 1.065 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 11.760 4.220 ;
        RECT 1.210 2.815 1.550 3.620 ;
        RECT 5.365 3.000 5.595 3.620 ;
        RECT 7.630 2.815 7.970 3.620 ;
        RECT 10.005 2.530 10.235 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 12.190 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.190 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 0.860 ;
        RECT 5.465 0.300 5.695 0.860 ;
        RECT 9.725 0.300 9.955 1.075 ;
        RECT 0.000 -0.300 11.760 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 2.580 0.530 3.380 ;
        RECT 3.160 3.095 4.560 3.325 ;
        RECT 0.190 2.350 3.160 2.580 ;
        RECT 0.190 0.530 0.530 2.350 ;
        RECT 4.320 1.455 4.560 3.095 ;
        RECT 6.665 2.580 6.895 3.380 ;
        RECT 8.605 2.625 8.835 3.250 ;
        RECT 4.810 2.350 7.970 2.580 ;
        RECT 8.605 2.395 9.755 2.625 ;
        RECT 7.630 2.145 7.970 2.350 ;
        RECT 7.630 1.805 9.285 2.145 ;
        RECT 9.525 2.020 9.755 2.395 ;
        RECT 4.320 1.225 6.530 1.455 ;
        RECT 4.320 0.760 4.560 1.225 ;
        RECT 3.410 0.530 4.560 0.760 ;
        RECT 7.630 0.530 7.970 1.805 ;
        RECT 9.525 1.790 10.750 2.020 ;
        RECT 9.525 1.555 9.755 1.790 ;
        RECT 8.605 1.325 9.755 1.555 ;
        RECT 8.605 0.735 8.835 1.325 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latsnq_1
MACRO gf180mcu_fd_sc_mcu7t5v0__latsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.320 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.965 1.790 3.270 2.120 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.293500 ;
    PORT
      LAYER Metal1 ;
        RECT 3.500 1.560 4.045 2.795 ;
        RECT 0.780 1.240 4.045 1.560 ;
    END
  END E
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.741500 ;
    PORT
      LAYER Metal1 ;
        RECT 5.040 1.800 7.380 2.120 ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.060800 ;
    PORT
      LAYER Metal1 ;
        RECT 10.640 2.340 11.100 3.380 ;
        RECT 10.640 2.110 11.660 2.340 ;
        RECT 11.300 1.380 11.660 2.110 ;
        RECT 10.640 1.130 11.660 1.380 ;
        RECT 10.640 0.555 11.100 1.130 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 12.320 4.220 ;
        RECT 1.365 3.000 1.595 3.620 ;
        RECT 5.365 3.000 5.595 3.620 ;
        RECT 7.630 2.815 7.970 3.620 ;
        RECT 9.525 2.570 9.755 3.620 ;
        RECT 11.665 2.570 11.895 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 12.750 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.750 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 0.860 ;
        RECT 5.465 0.300 5.695 0.860 ;
        RECT 9.525 0.300 9.755 0.895 ;
        RECT 11.765 0.300 11.995 0.895 ;
        RECT 0.000 -0.300 12.320 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 2.580 0.575 3.380 ;
        RECT 3.160 3.095 4.560 3.325 ;
        RECT 0.190 2.350 3.160 2.580 ;
        RECT 0.190 0.530 0.530 2.350 ;
        RECT 4.320 1.455 4.560 3.095 ;
        RECT 6.665 2.580 6.895 3.380 ;
        RECT 4.810 2.350 7.970 2.580 ;
        RECT 7.630 1.860 7.970 2.350 ;
        RECT 8.505 2.340 8.735 3.380 ;
        RECT 8.505 2.110 9.815 2.340 ;
        RECT 9.585 1.860 9.815 2.110 ;
        RECT 7.630 1.630 9.245 1.860 ;
        RECT 9.585 1.630 10.935 1.860 ;
        RECT 4.320 1.225 6.530 1.455 ;
        RECT 4.320 0.760 4.560 1.225 ;
        RECT 3.410 0.530 4.560 0.760 ;
        RECT 7.630 0.530 7.970 1.630 ;
        RECT 9.585 1.380 9.815 1.630 ;
        RECT 8.405 1.150 9.815 1.380 ;
        RECT 8.405 0.555 8.635 1.150 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latsnq_2
MACRO gf180mcu_fd_sc_mcu7t5v0__latsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.680 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.010 1.240 2.700 1.590 ;
        RECT 2.325 0.550 2.700 1.240 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.293500 ;
    PORT
      LAYER Metal1 ;
        RECT 3.490 2.120 4.045 2.795 ;
        RECT 0.780 1.820 4.045 2.120 ;
        RECT 2.950 1.270 3.210 1.820 ;
    END
  END E
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.040 1.800 7.390 2.120 ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.121600 ;
    PORT
      LAYER Metal1 ;
        RECT 11.860 2.340 12.220 3.380 ;
        RECT 13.965 2.340 14.460 3.380 ;
        RECT 11.860 2.110 15.000 2.340 ;
        RECT 14.670 1.390 15.000 2.110 ;
        RECT 11.825 1.160 15.000 1.390 ;
        RECT 11.825 0.545 12.055 1.160 ;
        RECT 14.065 0.545 14.295 1.160 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 15.680 4.220 ;
        RECT 1.365 3.000 1.595 3.620 ;
        RECT 5.590 2.815 5.930 3.620 ;
        RECT 7.630 2.815 7.970 3.620 ;
        RECT 8.565 2.570 8.795 3.620 ;
        RECT 10.755 2.570 10.985 3.620 ;
        RECT 12.945 2.570 13.175 3.620 ;
        RECT 14.985 2.570 15.215 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 16.110 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 16.110 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 1.115 ;
        RECT 5.410 0.300 5.750 1.065 ;
        RECT 8.465 0.300 8.695 0.885 ;
        RECT 10.705 0.300 10.935 0.885 ;
        RECT 12.945 0.300 13.175 0.885 ;
        RECT 15.185 0.300 15.415 0.885 ;
        RECT 0.000 -0.300 15.680 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 2.580 0.575 3.380 ;
        RECT 3.160 3.095 4.560 3.325 ;
        RECT 0.190 2.350 3.160 2.580 ;
        RECT 0.190 0.815 0.530 2.350 ;
        RECT 4.320 1.570 4.560 3.095 ;
        RECT 6.665 2.580 6.895 3.380 ;
        RECT 4.810 2.350 7.970 2.580 ;
        RECT 7.630 1.860 7.970 2.350 ;
        RECT 9.585 2.340 9.815 3.380 ;
        RECT 9.585 2.110 10.895 2.340 ;
        RECT 10.665 1.860 10.895 2.110 ;
        RECT 7.630 1.630 10.360 1.860 ;
        RECT 10.665 1.630 14.370 1.860 ;
        RECT 4.320 1.340 6.530 1.570 ;
        RECT 4.320 1.060 4.560 1.340 ;
        RECT 3.450 0.830 4.560 1.060 ;
        RECT 7.630 0.530 7.970 1.630 ;
        RECT 10.665 1.390 10.895 1.630 ;
        RECT 9.585 1.160 10.895 1.390 ;
        RECT 9.585 0.545 9.815 1.160 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latsnq_4
MACRO gf180mcu_fd_sc_mcu7t5v0__mux2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__mux2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.523500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.010 1.770 6.070 2.120 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.523500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.330 1.210 2.710 2.710 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.047000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.940 2.360 6.090 2.785 ;
        RECT 2.940 1.445 3.295 2.360 ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.130 0.650 0.575 3.270 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.280 4.220 ;
        RECT 1.365 2.760 1.595 3.620 ;
        RECT 5.310 3.105 5.650 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 7.710 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 0.865 ;
        RECT 5.465 0.300 5.695 0.880 ;
        RECT 0.000 -0.300 7.280 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.825 3.110 3.890 3.340 ;
        RECT 1.825 1.625 2.055 3.110 ;
        RECT 0.840 1.390 2.055 1.625 ;
        RECT 1.825 0.815 2.055 1.390 ;
        RECT 6.350 1.375 6.815 3.380 ;
        RECT 4.125 1.145 6.815 1.375 ;
        RECT 1.825 0.575 3.880 0.815 ;
        RECT 6.350 0.530 6.815 1.145 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__mux2_1
MACRO gf180mcu_fd_sc_mcu7t5v0__mux2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__mux2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.400 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.575 1.250 7.225 1.580 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.880 1.545 3.230 3.285 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.910 1.810 7.370 2.195 ;
        RECT 4.910 1.650 5.220 1.810 ;
        RECT 3.920 1.250 5.220 1.650 ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.121800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.250 0.540 1.650 3.380 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 8.400 4.220 ;
        RECT 0.295 2.530 0.525 3.620 ;
        RECT 2.385 2.530 2.615 3.620 ;
        RECT 6.590 2.965 6.930 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 8.830 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.830 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 0.835 ;
        RECT 2.485 0.300 2.715 0.835 ;
        RECT 6.645 0.300 6.875 0.835 ;
        RECT 0.000 -0.300 8.400 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.460 2.965 5.260 3.195 ;
        RECT 1.945 1.315 2.175 1.780 ;
        RECT 3.460 1.315 3.690 2.965 ;
        RECT 7.665 2.725 8.050 3.390 ;
        RECT 4.320 2.490 8.050 2.725 ;
        RECT 4.320 1.960 4.660 2.490 ;
        RECT 1.945 1.085 3.690 1.315 ;
        RECT 3.460 0.780 3.690 1.085 ;
        RECT 3.460 0.550 4.820 0.780 ;
        RECT 7.710 0.540 8.050 2.490 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__mux2_2
MACRO gf180mcu_fd_sc_mcu7t5v0__mux2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__mux2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.640 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.890 1.250 9.540 1.580 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.150 1.545 5.500 3.285 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.280 1.810 9.635 2.195 ;
        RECT 7.280 1.650 7.590 1.810 ;
        RECT 6.255 1.250 7.590 1.650 ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.304600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.250 2.120 1.705 3.380 ;
        RECT 3.490 2.120 3.945 3.380 ;
        RECT 1.250 1.800 3.945 2.120 ;
        RECT 1.250 0.540 1.705 1.800 ;
        RECT 3.490 0.540 3.945 1.800 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 10.640 4.220 ;
        RECT 0.350 2.530 0.580 3.620 ;
        RECT 2.490 2.530 2.720 3.620 ;
        RECT 4.680 2.530 4.910 3.620 ;
        RECT 8.885 2.955 9.225 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 11.070 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 11.070 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 0.300 0.530 0.835 ;
        RECT 2.540 0.300 2.770 0.835 ;
        RECT 4.780 0.300 5.010 0.835 ;
        RECT 8.940 0.300 9.170 0.835 ;
        RECT 0.000 -0.300 10.640 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 5.755 2.965 7.555 3.195 ;
        RECT 4.240 1.315 4.470 1.780 ;
        RECT 5.755 1.315 5.985 2.965 ;
        RECT 9.960 2.725 10.345 3.390 ;
        RECT 6.615 2.490 10.345 2.725 ;
        RECT 6.615 1.960 6.955 2.490 ;
        RECT 4.240 1.085 5.985 1.315 ;
        RECT 5.755 0.780 5.985 1.085 ;
        RECT 5.755 0.550 7.115 0.780 ;
        RECT 10.005 0.540 10.345 2.490 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__mux2_4
MACRO gf180mcu_fd_sc_mcu7t5v0__mux4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__mux4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.501500 ;
    PORT
      LAYER Metal1 ;
        RECT 15.250 1.750 16.940 2.120 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.501500 ;
    PORT
      LAYER Metal1 ;
        RECT 10.590 1.780 12.500 2.130 ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.501500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 0.970 1.010 2.950 ;
    END
  END I2
  PIN I3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.501500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.300 1.800 5.550 2.150 ;
        RECT 4.300 1.375 4.585 1.800 ;
    END
  END I3
  PIN S0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.504500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.185 2.120 2.415 2.465 ;
        RECT 2.185 1.800 3.495 2.120 ;
        RECT 3.200 1.240 3.495 1.800 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.003000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.070 2.150 9.300 2.465 ;
        RECT 7.960 1.770 9.300 2.150 ;
        RECT 7.960 1.165 8.300 1.770 ;
    END
  END S1
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.510400 ;
    PORT
      LAYER Metal1 ;
        RECT 5.990 1.570 6.380 2.855 ;
        RECT 5.650 0.600 6.380 1.570 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 17.920 4.220 ;
        RECT 0.245 2.685 0.475 3.620 ;
        RECT 4.845 2.845 5.185 3.620 ;
        RECT 11.670 2.845 12.015 3.620 ;
        RECT 15.955 2.815 16.295 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 18.350 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.130 ;
        RECT 4.850 0.300 5.080 1.160 ;
        RECT 11.630 0.300 11.860 1.145 ;
        RECT 16.110 0.300 16.340 1.145 ;
        RECT 0.000 -0.300 17.920 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.635 3.100 4.530 3.330 ;
        RECT 1.260 1.075 1.495 3.025 ;
        RECT 2.635 2.970 2.975 3.100 ;
        RECT 1.725 2.740 2.975 2.970 ;
        RECT 1.725 1.570 1.955 2.740 ;
        RECT 1.725 1.340 2.290 1.570 ;
        RECT 2.040 1.075 2.290 1.340 ;
        RECT 1.260 0.845 1.650 1.075 ;
        RECT 2.040 0.845 2.770 1.075 ;
        RECT 3.725 0.780 4.070 2.870 ;
        RECT 4.300 2.615 4.530 3.100 ;
        RECT 5.520 3.155 6.860 3.390 ;
        RECT 5.520 2.615 5.750 3.155 ;
        RECT 4.300 2.380 5.750 2.615 ;
        RECT 6.630 3.005 6.860 3.155 ;
        RECT 9.650 3.160 11.355 3.390 ;
        RECT 6.630 2.665 7.270 3.005 ;
        RECT 7.500 2.720 8.755 2.950 ;
        RECT 6.630 1.130 6.860 2.665 ;
        RECT 7.500 1.820 7.730 2.720 ;
        RECT 7.090 1.460 7.730 1.820 ;
        RECT 6.630 0.790 7.270 1.130 ;
        RECT 7.500 0.760 7.730 1.460 ;
        RECT 8.530 0.760 8.760 1.145 ;
        RECT 9.650 0.780 9.880 3.160 ;
        RECT 10.110 2.575 10.840 2.925 ;
        RECT 11.125 2.615 11.355 3.160 ;
        RECT 12.265 3.160 14.100 3.390 ;
        RECT 12.265 2.615 12.495 3.160 ;
        RECT 10.110 1.145 10.350 2.575 ;
        RECT 11.125 2.380 12.495 2.615 ;
        RECT 10.110 0.795 10.840 1.145 ;
        RECT 12.750 0.780 12.980 2.925 ;
        RECT 13.770 0.780 14.100 3.160 ;
        RECT 14.330 2.815 15.190 3.045 ;
        RECT 14.330 1.080 14.560 2.815 ;
        RECT 17.125 2.585 17.460 3.140 ;
        RECT 14.790 2.355 17.460 2.585 ;
        RECT 14.790 1.685 15.020 2.355 ;
        RECT 14.330 0.850 15.275 1.080 ;
        RECT 17.230 0.780 17.460 2.355 ;
        RECT 7.500 0.530 8.760 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__mux4_1
MACRO gf180mcu_fd_sc_mcu7t5v0__mux4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__mux4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.040 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.516500 ;
    PORT
      LAYER Metal1 ;
        RECT 16.485 1.780 18.175 2.120 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.516500 ;
    PORT
      LAYER Metal1 ;
        RECT 11.835 1.780 13.735 2.130 ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.618000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 0.970 1.010 2.950 ;
    END
  END I2
  PIN I3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.618000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.505 1.800 5.755 2.150 ;
        RECT 4.505 0.550 4.935 1.800 ;
    END
  END I3
  PIN S0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.651000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.255 1.800 3.700 2.250 ;
        RECT 3.300 1.240 3.700 1.800 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.033000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.165 2.150 10.535 3.320 ;
        RECT 9.170 1.770 10.535 2.150 ;
        RECT 9.170 1.305 9.535 1.770 ;
    END
  END S1
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.759200 ;
    PORT
      LAYER Metal1 ;
        RECT 6.230 0.600 6.600 2.855 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 19.040 4.220 ;
        RECT 0.245 2.575 0.475 3.620 ;
        RECT 5.010 2.845 5.350 3.620 ;
        RECT 7.405 2.570 7.635 3.620 ;
        RECT 12.905 2.845 13.250 3.620 ;
        RECT 17.190 2.815 17.530 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 19.470 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 19.470 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.130 ;
        RECT 5.165 0.300 5.395 1.160 ;
        RECT 7.405 0.300 7.635 1.160 ;
        RECT 12.865 0.300 13.095 1.145 ;
        RECT 17.345 0.300 17.575 1.145 ;
        RECT 0.000 -0.300 19.040 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.710 3.100 4.735 3.330 ;
        RECT 2.710 2.970 3.050 3.100 ;
        RECT 1.260 1.075 1.495 2.950 ;
        RECT 1.725 2.740 3.050 2.970 ;
        RECT 1.725 1.570 1.955 2.740 ;
        RECT 1.725 1.340 2.290 1.570 ;
        RECT 2.040 1.075 2.290 1.340 ;
        RECT 1.260 0.845 1.650 1.075 ;
        RECT 2.040 0.845 2.910 1.075 ;
        RECT 3.930 0.780 4.275 2.870 ;
        RECT 4.505 2.615 4.735 3.100 ;
        RECT 5.670 3.155 7.095 3.390 ;
        RECT 5.670 2.615 5.900 3.155 ;
        RECT 4.505 2.380 5.900 2.615 ;
        RECT 6.865 2.275 7.095 3.155 ;
        RECT 10.885 3.160 12.590 3.390 ;
        RECT 7.865 2.665 8.480 3.005 ;
        RECT 8.710 2.720 9.880 2.950 ;
        RECT 7.865 2.275 8.095 2.665 ;
        RECT 6.865 2.045 8.095 2.275 ;
        RECT 7.865 1.130 8.095 2.045 ;
        RECT 8.710 1.820 8.940 2.720 ;
        RECT 8.325 1.460 8.940 1.820 ;
        RECT 7.865 0.790 8.480 1.130 ;
        RECT 8.710 1.075 8.940 1.460 ;
        RECT 8.710 0.845 9.950 1.075 ;
        RECT 10.885 0.780 11.115 3.160 ;
        RECT 11.345 2.575 12.075 2.925 ;
        RECT 12.360 2.615 12.590 3.160 ;
        RECT 13.500 3.160 15.335 3.390 ;
        RECT 13.500 2.615 13.730 3.160 ;
        RECT 11.345 1.145 11.595 2.575 ;
        RECT 12.360 2.380 13.730 2.615 ;
        RECT 11.345 0.795 12.075 1.145 ;
        RECT 13.985 0.780 14.215 2.925 ;
        RECT 15.005 0.780 15.335 3.160 ;
        RECT 15.565 2.815 16.425 3.045 ;
        RECT 15.565 1.080 15.795 2.815 ;
        RECT 18.360 2.585 18.695 3.140 ;
        RECT 16.025 2.355 18.695 2.585 ;
        RECT 16.025 1.675 16.255 2.355 ;
        RECT 15.565 0.850 16.510 1.080 ;
        RECT 18.465 0.780 18.695 2.355 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__mux4_2
MACRO gf180mcu_fd_sc_mcu7t5v0__mux4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__mux4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.516500 ;
    PORT
      LAYER Metal1 ;
        RECT 18.725 1.780 20.415 2.120 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.516500 ;
    PORT
      LAYER Metal1 ;
        RECT 14.075 1.780 15.975 2.130 ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.618000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 1.025 1.010 2.835 ;
    END
  END I2
  PIN I3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.618000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.505 1.800 5.755 2.150 ;
        RECT 4.505 0.550 4.935 1.800 ;
    END
  END I3
  PIN S0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.651000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.255 1.800 3.700 2.250 ;
        RECT 3.300 1.240 3.700 1.800 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.033000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.405 2.150 12.775 3.320 ;
        RECT 11.410 1.770 12.775 2.150 ;
        RECT 11.410 1.305 11.775 1.770 ;
    END
  END S1
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.206400 ;
    PORT
      LAYER Metal1 ;
        RECT 6.230 2.150 6.615 2.925 ;
        RECT 8.425 2.150 8.840 2.925 ;
        RECT 6.230 1.800 8.840 2.150 ;
        RECT 6.230 0.600 6.600 1.800 ;
        RECT 8.425 0.600 8.840 1.800 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 21.280 4.220 ;
        RECT 0.245 2.575 0.475 3.620 ;
        RECT 5.120 2.845 5.460 3.620 ;
        RECT 7.350 2.845 7.690 3.620 ;
        RECT 9.530 2.845 9.870 3.620 ;
        RECT 15.145 2.845 15.490 3.620 ;
        RECT 19.430 2.815 19.770 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 21.710 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.710 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.130 ;
        RECT 5.165 0.300 5.395 1.160 ;
        RECT 7.405 0.300 7.635 1.160 ;
        RECT 9.645 0.300 9.875 1.160 ;
        RECT 15.105 0.300 15.335 1.145 ;
        RECT 19.585 0.300 19.815 1.145 ;
        RECT 0.000 -0.300 21.280 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.710 3.100 4.735 3.330 ;
        RECT 2.710 2.970 3.050 3.100 ;
        RECT 1.260 1.075 1.495 2.950 ;
        RECT 1.725 2.740 3.050 2.970 ;
        RECT 1.725 1.570 1.955 2.740 ;
        RECT 1.725 1.340 2.290 1.570 ;
        RECT 2.040 1.075 2.290 1.340 ;
        RECT 1.260 0.845 1.650 1.075 ;
        RECT 2.040 0.845 2.910 1.075 ;
        RECT 3.930 0.780 4.275 2.870 ;
        RECT 4.505 2.615 4.735 3.100 ;
        RECT 5.755 3.160 7.120 3.390 ;
        RECT 5.755 2.615 5.985 3.160 ;
        RECT 4.505 2.380 5.985 2.615 ;
        RECT 6.890 2.615 7.120 3.160 ;
        RECT 7.920 3.155 9.300 3.390 ;
        RECT 7.920 2.615 8.150 3.155 ;
        RECT 6.890 2.380 8.150 2.615 ;
        RECT 9.070 2.615 9.300 3.155 ;
        RECT 13.125 3.160 14.830 3.390 ;
        RECT 10.490 2.615 10.720 3.005 ;
        RECT 9.070 2.380 10.720 2.615 ;
        RECT 10.950 2.720 12.120 2.950 ;
        RECT 10.105 1.130 10.335 2.380 ;
        RECT 10.950 1.820 11.180 2.720 ;
        RECT 10.565 1.460 11.180 1.820 ;
        RECT 10.105 0.790 10.720 1.130 ;
        RECT 10.950 1.075 11.180 1.460 ;
        RECT 10.950 0.845 12.190 1.075 ;
        RECT 13.125 0.780 13.355 3.160 ;
        RECT 13.585 2.575 14.315 2.925 ;
        RECT 14.600 2.615 14.830 3.160 ;
        RECT 15.740 3.160 17.575 3.390 ;
        RECT 15.740 2.615 15.970 3.160 ;
        RECT 13.585 1.145 13.835 2.575 ;
        RECT 14.600 2.380 15.970 2.615 ;
        RECT 13.585 0.795 14.315 1.145 ;
        RECT 16.225 0.780 16.455 2.925 ;
        RECT 17.245 0.780 17.575 3.160 ;
        RECT 17.805 2.815 18.665 3.045 ;
        RECT 17.805 1.080 18.035 2.815 ;
        RECT 20.600 2.585 20.935 3.140 ;
        RECT 18.265 2.355 20.935 2.585 ;
        RECT 18.265 1.675 18.495 2.355 ;
        RECT 17.805 0.850 18.750 1.080 ;
        RECT 20.705 0.780 20.935 2.355 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__mux4_4
MACRO gf180mcu_fd_sc_mcu7t5v0__nand2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nand2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.800 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.057000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.240 1.440 2.055 1.820 ;
        RECT 1.240 0.555 1.605 1.440 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.057000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 1.060 1.000 2.190 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.948400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 2.300 1.500 3.380 ;
        RECT 1.270 2.070 2.680 2.300 ;
        RECT 2.290 0.530 2.680 2.070 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 2.800 4.220 ;
        RECT 0.250 2.530 0.480 3.620 ;
        RECT 2.290 2.530 2.520 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 3.230 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 3.230 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 0.300 0.480 0.805 ;
        RECT 0.000 -0.300 2.800 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nand2_1
MACRO gf180mcu_fd_sc_mcu7t5v0__nand2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nand2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.040 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.114000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.620 1.240 3.160 1.560 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.114000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.620 1.800 4.030 2.120 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.601600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.220 2.680 1.580 3.380 ;
        RECT 3.305 2.680 3.535 3.380 ;
        RECT 1.220 2.360 4.490 2.680 ;
        RECT 4.260 1.535 4.490 2.360 ;
        RECT 3.460 1.265 4.490 1.535 ;
        RECT 3.460 1.000 3.820 1.265 ;
        RECT 2.150 0.680 3.820 1.000 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.040 4.220 ;
        RECT 0.245 2.640 0.475 3.620 ;
        RECT 2.285 3.085 2.515 3.620 ;
        RECT 4.325 3.085 4.555 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 5.470 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 5.470 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 0.905 ;
        RECT 4.260 0.300 4.620 0.635 ;
        RECT 0.000 -0.300 5.040 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nand2_2
MACRO gf180mcu_fd_sc_mcu7t5v0__nand2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nand2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.960 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.228000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 1.800 7.175 2.130 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.228000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.405 1.825 8.110 2.095 ;
        RECT 7.405 1.570 7.635 1.825 ;
        RECT 0.610 1.325 7.635 1.570 ;
        RECT 0.610 1.240 3.545 1.325 ;
        RECT 5.265 1.240 7.635 1.325 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.240100 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 2.680 1.495 3.390 ;
        RECT 3.305 2.680 3.535 3.390 ;
        RECT 5.345 2.680 5.575 3.390 ;
        RECT 7.385 2.680 7.615 3.390 ;
        RECT 1.265 2.360 8.570 2.680 ;
        RECT 8.340 1.575 8.570 2.360 ;
        RECT 7.885 1.345 8.570 1.575 ;
        RECT 3.775 1.010 5.035 1.095 ;
        RECT 7.885 1.010 8.115 1.345 ;
        RECT 2.140 0.865 8.115 1.010 ;
        RECT 2.140 0.680 4.005 0.865 ;
        RECT 4.805 0.680 8.115 0.865 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 8.960 4.220 ;
        RECT 0.245 2.640 0.475 3.620 ;
        RECT 2.285 2.930 2.515 3.620 ;
        RECT 4.325 2.930 4.555 3.620 ;
        RECT 6.365 2.930 6.595 3.620 ;
        RECT 8.405 2.930 8.635 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 9.390 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.390 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.325 0.300 0.555 0.905 ;
        RECT 4.235 0.300 4.575 0.635 ;
        RECT 8.350 0.300 8.690 0.635 ;
        RECT 0.000 -0.300 8.960 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nand2_4
MACRO gf180mcu_fd_sc_mcu7t5v0__nand3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nand3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.920 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.984500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.900 0.550 3.210 1.960 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.984500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.780 0.550 2.140 1.960 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.984500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.120 1.760 1.065 2.150 ;
        RECT 0.660 1.055 1.065 1.760 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.306400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 2.780 1.630 3.380 ;
        RECT 3.380 2.780 3.670 3.380 ;
        RECT 1.400 2.360 3.670 2.780 ;
        RECT 3.440 0.655 3.670 2.360 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 3.920 4.220 ;
        RECT 0.380 2.530 0.610 3.620 ;
        RECT 2.365 3.130 2.705 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 4.350 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.350 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.380 0.300 0.610 0.805 ;
        RECT 0.000 -0.300 3.920 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nand3_1
MACRO gf180mcu_fd_sc_mcu7t5v0__nand3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nand3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.969000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.950 1.265 4.200 1.555 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.969000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.770 1.785 5.050 2.020 ;
        RECT 4.530 1.535 5.050 1.785 ;
        RECT 4.530 1.260 6.245 1.535 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.969000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 2.250 6.175 2.485 ;
        RECT 1.265 2.150 1.540 2.250 ;
        RECT 0.780 1.770 1.540 2.150 ;
        RECT 5.690 2.150 6.175 2.250 ;
        RECT 5.690 1.785 6.670 2.150 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.963000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.130 2.715 5.725 2.950 ;
        RECT 0.130 1.100 0.430 2.715 ;
        RECT 0.130 0.975 1.370 1.100 ;
        RECT 0.130 0.865 3.995 0.975 ;
        RECT 1.040 0.705 3.995 0.865 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.280 4.220 ;
        RECT 0.265 3.180 0.495 3.620 ;
        RECT 2.305 3.180 2.535 3.620 ;
        RECT 4.345 3.180 4.575 3.620 ;
        RECT 6.385 2.640 6.615 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 7.710 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 0.300 0.690 0.635 ;
        RECT 6.385 0.300 6.615 0.900 ;
        RECT 0.000 -0.300 7.280 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nand3_2
MACRO gf180mcu_fd_sc_mcu7t5v0__nand3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nand3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.938000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.050 1.790 12.670 2.130 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.938000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 1.790 8.530 2.150 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.938000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.710 1.330 7.540 1.560 ;
        RECT 3.450 1.210 5.660 1.330 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.801400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.210 2.755 1.550 3.360 ;
        RECT 3.350 2.755 3.690 3.360 ;
        RECT 5.490 2.755 5.830 3.360 ;
        RECT 7.630 2.755 7.970 3.360 ;
        RECT 9.990 2.755 10.330 3.360 ;
        RECT 12.660 2.755 13.350 3.360 ;
        RECT 1.210 2.380 13.350 2.755 ;
        RECT 12.970 1.220 13.350 2.380 ;
        RECT 9.680 0.990 13.350 1.220 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 14.560 4.220 ;
        RECT 0.245 2.760 0.475 3.620 ;
        RECT 2.285 2.985 2.515 3.620 ;
        RECT 4.425 2.985 4.655 3.620 ;
        RECT 6.565 2.985 6.795 3.620 ;
        RECT 8.705 2.985 8.935 3.620 ;
        RECT 11.285 2.985 11.515 3.620 ;
        RECT 13.965 2.760 14.195 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 14.990 4.350 ;
        RECT -0.430 1.760 9.610 1.885 ;
        RECT 13.390 1.760 14.990 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 9.610 1.760 13.390 1.885 ;
        RECT -0.430 -0.430 14.990 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.320 0.300 2.680 0.635 ;
        RECT 6.600 0.300 6.960 0.635 ;
        RECT 0.000 -0.300 14.560 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.180 0.865 3.175 1.095 ;
        RECT 2.945 0.760 3.175 0.865 ;
        RECT 6.135 0.865 7.980 1.100 ;
        RECT 6.135 0.760 6.365 0.865 ;
        RECT 2.945 0.530 6.365 0.760 ;
        RECT 7.750 0.760 7.980 0.865 ;
        RECT 7.750 0.530 14.360 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__nand3_4
MACRO gf180mcu_fd_sc_mcu7t5v0__nand4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nand4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.040 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.914500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.020 1.210 4.370 2.190 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.914500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.900 0.610 3.240 2.190 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.914500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 0.610 2.140 2.190 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.914500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.660 1.890 1.400 2.190 ;
        RECT 0.660 1.210 1.020 1.890 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.239600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.260 2.945 1.650 3.390 ;
        RECT 3.460 2.950 3.770 3.390 ;
        RECT 3.460 2.945 4.910 2.950 ;
        RECT 1.260 2.715 4.910 2.945 ;
        RECT 4.600 0.980 4.910 2.715 ;
        RECT 3.775 0.530 4.910 0.980 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.040 4.220 ;
        RECT 0.400 3.180 0.630 3.620 ;
        RECT 2.440 3.180 2.670 3.620 ;
        RECT 4.480 3.180 4.710 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 5.470 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 5.470 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 0.300 0.630 0.980 ;
        RECT 0.000 -0.300 5.040 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nand4_1
MACRO gf180mcu_fd_sc_mcu7t5v0__nand4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nand4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.960 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.829000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.610 1.820 2.580 2.100 ;
        RECT 2.350 1.675 2.580 1.820 ;
        RECT 2.350 1.445 4.030 1.675 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.829000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.810 1.905 5.775 2.135 ;
        RECT 4.455 1.750 5.775 1.905 ;
        RECT 5.500 1.695 5.775 1.750 ;
        RECT 5.500 1.465 6.150 1.695 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.829000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.610 1.215 2.095 1.590 ;
        RECT 6.810 1.220 7.190 1.555 ;
        RECT 4.080 1.215 7.190 1.220 ;
        RECT 0.610 1.210 7.190 1.215 ;
        RECT 1.755 0.990 7.190 1.210 ;
        RECT 1.755 0.985 4.130 0.990 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.829000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.690 2.365 6.660 2.595 ;
        RECT 0.690 2.340 1.845 2.365 ;
        RECT 6.380 2.260 6.660 2.365 ;
        RECT 6.380 1.825 8.190 2.260 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.488200 ;
    PORT
      LAYER Metal1 ;
        RECT 0.180 3.055 0.980 3.310 ;
        RECT 1.810 3.055 3.020 3.310 ;
        RECT 3.935 3.055 4.900 3.310 ;
        RECT 6.055 3.055 7.140 3.310 ;
        RECT 0.180 2.825 7.140 3.055 ;
        RECT 6.910 2.760 7.140 2.825 ;
        RECT 8.405 2.760 8.815 3.390 ;
        RECT 6.910 2.525 8.815 2.760 ;
        RECT 8.495 1.535 8.815 2.525 ;
        RECT 7.425 1.265 8.815 1.535 ;
        RECT 7.425 0.760 7.695 1.265 ;
        RECT 4.180 0.530 7.695 0.760 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 8.960 4.220 ;
        RECT 1.210 3.285 1.550 3.620 ;
        RECT 3.250 3.285 3.590 3.620 ;
        RECT 5.290 3.285 5.630 3.620 ;
        RECT 7.385 3.000 7.615 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 9.390 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.390 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 0.830 ;
        RECT 8.405 0.300 8.635 0.830 ;
        RECT 0.000 -0.300 8.960 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nand4_2
MACRO gf180mcu_fd_sc_mcu7t5v0__nand4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nand4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.658000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.950 1.535 16.155 1.680 ;
        RECT 8.450 1.450 16.155 1.535 ;
        RECT 8.450 1.265 10.300 1.450 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.658000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.450 1.910 17.270 2.150 ;
        RECT 8.450 1.825 9.470 1.910 ;
        RECT 16.385 1.750 17.270 1.910 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.658000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.620 1.825 8.200 2.095 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.658000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.730 1.325 7.180 1.555 ;
        RECT 3.345 1.210 5.510 1.325 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.179600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 2.655 1.495 3.310 ;
        RECT 3.305 2.655 3.535 3.310 ;
        RECT 5.345 2.655 5.575 3.310 ;
        RECT 7.385 2.655 7.615 3.310 ;
        RECT 9.425 2.655 9.655 3.310 ;
        RECT 11.905 2.655 12.135 3.310 ;
        RECT 13.945 2.655 14.175 3.310 ;
        RECT 16.425 2.655 16.655 3.310 ;
        RECT 1.265 2.380 17.775 2.655 ;
        RECT 17.505 1.220 17.775 2.380 ;
        RECT 10.600 0.990 17.775 1.220 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 17.920 4.220 ;
        RECT 0.245 2.840 0.475 3.620 ;
        RECT 2.285 2.935 2.515 3.620 ;
        RECT 4.325 2.935 4.555 3.620 ;
        RECT 6.365 2.935 6.595 3.620 ;
        RECT 8.405 2.935 8.635 3.620 ;
        RECT 10.885 2.935 11.115 3.620 ;
        RECT 12.925 2.935 13.155 3.620 ;
        RECT 15.405 2.935 15.635 3.620 ;
        RECT 17.445 2.935 17.675 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 18.350 4.350 ;
        RECT -0.430 1.760 10.230 1.885 ;
        RECT 15.850 1.760 18.350 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 10.230 1.760 15.850 1.885 ;
        RECT -0.430 -0.430 18.350 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.220 0.300 2.580 0.635 ;
        RECT 6.300 0.300 6.660 0.635 ;
        RECT 0.000 -0.300 17.920 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.180 0.980 3.040 1.095 ;
        RECT 5.840 0.980 7.635 1.095 ;
        RECT 0.180 0.865 7.635 0.980 ;
        RECT 2.810 0.690 6.070 0.865 ;
        RECT 7.405 0.760 7.635 0.865 ;
        RECT 7.405 0.530 17.730 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__nand4_4
MACRO gf180mcu_fd_sc_mcu7t5v0__nor2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.949000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.825 1.790 2.855 2.130 ;
        RECT 1.825 0.600 2.130 1.790 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.949000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 1.180 1.010 3.320 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.830600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.385 2.680 2.665 3.380 ;
        RECT 1.240 2.360 2.665 2.680 ;
        RECT 1.240 0.600 1.595 2.360 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 3.360 4.220 ;
        RECT 0.245 2.530 0.475 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 3.790 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 3.790 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 0.945 ;
        RECT 2.485 0.300 2.715 1.090 ;
        RECT 0.000 -0.300 3.360 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nor2_1
MACRO gf180mcu_fd_sc_mcu7t5v0__nor2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.898000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.480 1.770 3.220 2.150 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.898000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.810 2.380 3.780 2.700 ;
        RECT 0.810 1.580 1.060 2.380 ;
        RECT 3.480 2.150 3.780 2.380 ;
        RECT 3.480 1.770 4.390 2.150 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.283000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.390 3.140 4.325 3.370 ;
        RECT 4.095 3.035 4.325 3.140 ;
        RECT 4.095 2.800 4.895 3.035 ;
        RECT 4.625 1.320 4.895 2.800 ;
        RECT 1.365 1.050 4.895 1.320 ;
        RECT 1.365 0.530 1.595 1.050 ;
        RECT 3.605 0.530 3.835 1.050 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.600 4.220 ;
        RECT 0.295 2.625 0.525 3.620 ;
        RECT 4.610 3.285 4.970 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 6.030 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.180 0.300 0.540 0.820 ;
        RECT 2.420 0.300 2.780 0.820 ;
        RECT 4.660 0.300 5.020 0.820 ;
        RECT 0.000 -0.300 5.600 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nor2_2
MACRO gf180mcu_fd_sc_mcu7t5v0__nor2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.796000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.650 1.800 8.415 2.120 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.796000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.060 1.560 9.420 2.255 ;
        RECT 0.795 1.325 9.420 1.560 ;
        RECT 8.040 1.220 9.420 1.325 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.932000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.485 2.700 2.715 3.380 ;
        RECT 6.965 2.700 7.195 3.380 ;
        RECT 1.170 2.585 3.870 2.700 ;
        RECT 5.650 2.585 7.195 2.700 ;
        RECT 0.130 2.350 7.195 2.585 ;
        RECT 0.130 1.095 0.430 2.350 ;
        RECT 0.130 0.865 7.730 1.095 ;
        RECT 1.365 0.530 1.595 0.865 ;
        RECT 3.605 0.530 3.835 0.865 ;
        RECT 5.845 0.530 6.075 0.865 ;
        RECT 7.500 0.760 7.730 0.865 ;
        RECT 7.500 0.530 8.410 0.760 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 10.080 4.220 ;
        RECT 0.240 2.815 0.580 3.620 ;
        RECT 4.670 2.815 5.010 3.620 ;
        RECT 9.100 2.815 9.440 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 10.510 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.180 0.300 0.540 0.635 ;
        RECT 2.430 0.300 2.770 0.635 ;
        RECT 4.670 0.300 5.010 0.635 ;
        RECT 6.910 0.300 7.250 0.635 ;
        RECT 9.140 0.300 9.500 0.635 ;
        RECT 0.000 -0.300 10.080 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nor2_4
MACRO gf180mcu_fd_sc_mcu7t5v0__nor3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.889000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.910 1.575 3.250 3.390 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.889000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.790 1.575 2.130 3.390 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.889000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.220 2.190 1.560 3.390 ;
        RECT 0.490 1.760 1.560 2.190 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.983200 ;
    PORT
      LAYER Metal1 ;
        RECT 3.490 1.285 3.890 3.390 ;
        RECT 1.310 1.050 3.890 1.285 ;
        RECT 1.310 0.695 1.650 1.050 ;
        RECT 3.550 0.695 3.890 1.050 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 4.480 4.220 ;
        RECT 0.345 2.530 0.575 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 4.910 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 0.820 ;
        RECT 2.430 0.300 2.770 0.820 ;
        RECT 0.000 -0.300 4.480 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nor3_1
MACRO gf180mcu_fd_sc_mcu7t5v0__nor3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.955 1.825 4.390 2.095 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.935 1.770 2.710 2.095 ;
        RECT 2.385 1.590 2.710 1.770 ;
        RECT 4.625 1.770 5.650 2.150 ;
        RECT 4.625 1.590 4.895 1.770 ;
        RECT 2.385 1.360 4.895 1.590 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.305 2.380 6.630 2.655 ;
        RECT 1.305 1.665 1.580 2.380 ;
        RECT 6.250 1.730 6.630 2.380 ;
        RECT 0.705 1.390 1.580 1.665 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.649200 ;
    PORT
      LAYER Metal1 ;
        RECT 0.825 2.940 3.840 3.235 ;
        RECT 0.825 2.250 1.055 2.940 ;
        RECT 0.145 2.020 1.055 2.250 ;
        RECT 0.145 1.115 0.420 2.020 ;
        RECT 0.145 0.885 7.250 1.115 ;
        RECT 0.145 0.530 0.530 0.885 ;
        RECT 1.890 0.530 3.310 0.885 ;
        RECT 4.130 0.530 5.550 0.885 ;
        RECT 6.905 0.530 7.250 0.885 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.840 4.220 ;
        RECT 0.345 2.590 0.575 3.620 ;
        RECT 6.865 2.630 7.095 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 8.270 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.300 0.300 1.660 0.655 ;
        RECT 3.540 0.300 3.900 0.655 ;
        RECT 5.780 0.300 6.140 0.655 ;
        RECT 0.000 -0.300 7.840 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nor3_2
MACRO gf180mcu_fd_sc_mcu7t5v0__nor3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.556000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.550 1.640 9.960 2.850 ;
        RECT 9.550 1.410 12.180 1.640 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.556000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.405 1.870 9.030 2.150 ;
        RECT 0.405 1.750 1.570 1.870 ;
        RECT 7.970 1.750 9.030 1.870 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.556000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.790 1.410 7.735 1.640 ;
        RECT 3.470 1.010 3.910 1.410 ;
        RECT 5.700 1.010 6.150 1.410 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.963600 ;
    PORT
      LAYER Metal1 ;
        RECT 10.190 2.110 10.555 2.910 ;
        RECT 12.460 2.110 12.850 2.910 ;
        RECT 10.190 1.875 12.850 2.110 ;
        RECT 12.420 1.180 12.850 1.875 ;
        RECT 1.255 0.945 3.230 1.180 ;
        RECT 1.255 0.530 1.650 0.945 ;
        RECT 3.000 0.760 3.230 0.945 ;
        RECT 4.210 0.945 5.470 1.180 ;
        RECT 4.210 0.760 4.440 0.945 ;
        RECT 3.000 0.530 4.440 0.760 ;
        RECT 5.240 0.760 5.470 0.945 ;
        RECT 6.450 0.945 12.850 1.180 ;
        RECT 6.450 0.760 6.680 0.945 ;
        RECT 5.240 0.530 6.680 0.760 ;
        RECT 7.950 0.530 8.820 0.945 ;
        RECT 9.720 0.530 11.160 0.945 ;
        RECT 12.460 0.530 12.850 0.945 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 14.560 4.220 ;
        RECT 2.385 3.155 2.615 3.620 ;
        RECT 6.865 3.155 7.095 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 14.990 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 0.655 ;
        RECT 2.430 0.300 2.770 0.655 ;
        RECT 4.670 0.300 5.010 0.655 ;
        RECT 6.910 0.300 7.250 0.655 ;
        RECT 9.150 0.300 9.490 0.655 ;
        RECT 11.390 0.300 11.730 0.655 ;
        RECT 13.630 0.300 13.970 0.655 ;
        RECT 0.000 -0.300 14.560 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 2.800 0.475 3.380 ;
        RECT 4.625 2.800 4.855 3.380 ;
        RECT 7.990 3.160 13.815 3.390 ;
        RECT 7.990 2.800 8.220 3.160 ;
        RECT 0.245 2.570 8.220 2.800 ;
        RECT 11.345 2.530 11.575 3.160 ;
        RECT 13.585 2.530 13.815 3.160 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__nor3_4
MACRO gf180mcu_fd_sc_mcu7t5v0__nor4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.826000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.030 1.685 4.370 3.380 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.826000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.910 1.685 3.250 3.380 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.826000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.790 1.685 2.130 3.380 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.826000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.220 2.195 1.560 3.380 ;
        RECT 0.585 1.685 1.560 2.195 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.911200 ;
    PORT
      LAYER Metal1 ;
        RECT 4.610 2.380 4.905 3.380 ;
        RECT 4.610 1.305 4.910 2.380 ;
        RECT 1.255 1.070 4.910 1.305 ;
        RECT 1.255 0.530 1.650 1.070 ;
        RECT 3.505 0.530 3.890 1.070 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.600 4.220 ;
        RECT 0.345 2.530 0.575 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 6.030 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 0.840 ;
        RECT 2.485 0.300 2.715 0.840 ;
        RECT 4.725 0.300 4.955 0.840 ;
        RECT 0.000 -0.300 5.600 0.300 ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nor4_1
MACRO gf180mcu_fd_sc_mcu7t5v0__nor4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.652000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.835 1.560 8.745 1.695 ;
        RECT 6.835 1.465 9.630 1.560 ;
        RECT 8.470 1.240 9.630 1.465 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.652000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.690 1.930 9.630 2.160 ;
        RECT 5.690 1.750 6.605 1.930 ;
        RECT 8.975 1.800 9.630 1.930 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.652000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.385 1.930 4.615 2.160 ;
        RECT 0.385 1.825 1.275 1.930 ;
        RECT 3.450 1.825 4.615 1.930 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.652000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.505 1.565 3.220 1.695 ;
        RECT 0.385 1.465 3.220 1.565 ;
        RECT 0.385 1.265 1.735 1.465 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.631000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.130 2.390 7.790 2.665 ;
        RECT 5.130 1.235 5.460 2.390 ;
        RECT 1.975 1.005 3.235 1.235 ;
        RECT 1.975 0.975 2.205 1.005 ;
        RECT 1.170 0.530 2.205 0.975 ;
        RECT 3.005 0.975 3.235 1.005 ;
        RECT 4.395 1.005 5.655 1.235 ;
        RECT 4.395 0.975 4.625 1.005 ;
        RECT 3.005 0.530 4.625 0.975 ;
        RECT 5.425 0.975 5.655 1.005 ;
        RECT 6.815 1.005 8.145 1.235 ;
        RECT 6.815 0.975 7.045 1.005 ;
        RECT 5.425 0.530 7.045 0.975 ;
        RECT 7.845 0.975 8.145 1.005 ;
        RECT 7.845 0.530 8.950 0.975 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 10.080 4.220 ;
        RECT 2.440 2.935 2.670 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 10.510 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.195 0.300 0.535 0.775 ;
        RECT 2.435 0.300 2.775 0.775 ;
        RECT 4.855 0.300 5.195 0.775 ;
        RECT 7.275 0.300 7.615 0.775 ;
        RECT 9.515 0.300 9.855 0.775 ;
        RECT 0.000 -0.300 10.080 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.350 2.625 0.580 3.380 ;
        RECT 9.470 3.195 9.700 3.380 ;
        RECT 4.385 2.965 9.700 3.195 ;
        RECT 4.385 2.625 4.615 2.965 ;
        RECT 0.350 2.390 4.615 2.625 ;
        RECT 9.470 2.530 9.700 2.965 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__nor4_2
MACRO gf180mcu_fd_sc_mcu7t5v0__nor4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.720 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.294000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.855 1.535 18.890 1.680 ;
        RECT 11.855 1.450 20.110 1.535 ;
        RECT 13.545 1.170 13.890 1.450 ;
        RECT 16.325 1.170 16.685 1.450 ;
        RECT 18.660 1.265 20.110 1.450 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.294000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.510 1.910 20.110 2.150 ;
        RECT 10.510 1.770 11.625 1.910 ;
        RECT 19.140 1.770 20.110 1.910 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.294000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.610 1.910 9.395 2.150 ;
        RECT 0.610 1.820 1.295 1.910 ;
        RECT 8.460 1.730 9.395 1.910 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.294000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.540 1.535 8.210 1.680 ;
        RECT 0.610 1.450 8.210 1.535 ;
        RECT 0.610 1.265 1.760 1.450 ;
        RECT 3.510 1.170 3.850 1.450 ;
        RECT 6.240 1.170 6.585 1.450 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.830400 ;
    PORT
      LAYER Metal1 ;
        RECT 12.570 2.665 12.910 2.840 ;
        RECT 9.660 2.655 12.910 2.665 ;
        RECT 17.215 2.655 18.070 2.835 ;
        RECT 9.660 2.380 18.070 2.655 ;
        RECT 9.660 1.520 10.240 2.380 ;
        RECT 9.660 1.480 11.070 1.520 ;
        RECT 8.535 1.220 11.070 1.480 ;
        RECT 2.020 0.990 3.280 1.220 ;
        RECT 2.020 0.975 2.250 0.990 ;
        RECT 1.170 0.530 2.250 0.975 ;
        RECT 3.050 0.920 3.280 0.990 ;
        RECT 4.440 0.990 5.700 1.220 ;
        RECT 4.440 0.920 4.670 0.990 ;
        RECT 3.050 0.530 4.670 0.920 ;
        RECT 5.470 0.920 5.700 0.990 ;
        RECT 6.860 0.990 8.120 1.220 ;
        RECT 6.860 0.920 7.090 0.990 ;
        RECT 5.470 0.530 7.090 0.920 ;
        RECT 7.890 0.975 8.120 0.990 ;
        RECT 8.535 0.990 13.240 1.220 ;
        RECT 8.535 0.975 9.510 0.990 ;
        RECT 7.890 0.530 9.510 0.975 ;
        RECT 10.405 0.530 12.210 0.990 ;
        RECT 13.010 0.920 13.240 0.990 ;
        RECT 14.570 0.990 15.830 1.220 ;
        RECT 14.570 0.920 14.800 0.990 ;
        RECT 13.010 0.530 14.800 0.920 ;
        RECT 15.600 0.920 15.830 0.990 ;
        RECT 17.160 0.990 18.430 1.220 ;
        RECT 17.160 0.920 17.390 0.990 ;
        RECT 15.600 0.530 17.390 0.920 ;
        RECT 18.200 0.975 18.430 0.990 ;
        RECT 18.200 0.530 19.550 0.975 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 20.720 4.220 ;
        RECT 2.485 2.950 2.715 3.620 ;
        RECT 7.325 2.950 7.555 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 21.150 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.150 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.240 0.300 0.580 0.760 ;
        RECT 2.480 0.300 2.820 0.760 ;
        RECT 4.900 0.300 5.240 0.760 ;
        RECT 7.320 0.300 7.660 0.760 ;
        RECT 9.835 0.300 10.175 0.760 ;
        RECT 12.440 0.300 12.780 0.760 ;
        RECT 15.030 0.300 15.370 0.760 ;
        RECT 17.630 0.300 17.970 0.760 ;
        RECT 20.140 0.300 20.480 0.760 ;
        RECT 0.000 -0.300 20.720 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.395 2.650 0.625 3.380 ;
        RECT 4.905 2.650 5.135 3.390 ;
        RECT 8.510 3.150 20.380 3.385 ;
        RECT 8.510 2.650 8.740 3.150 ;
        RECT 14.890 2.945 15.230 3.150 ;
        RECT 0.395 2.415 8.740 2.650 ;
        RECT 20.040 2.530 20.380 3.150 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__nor4_4
MACRO gf180mcu_fd_sc_mcu7t5v0__oai21_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai21_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.825 0.550 2.160 2.320 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 0.550 1.000 2.230 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.057000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.375 1.900 4.350 2.150 ;
        RECT 2.945 1.600 4.350 1.900 ;
        RECT 2.945 0.550 3.280 1.600 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.230 2.590 2.615 2.930 ;
        RECT 1.230 0.550 1.595 2.590 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 4.480 4.220 ;
        RECT 0.295 2.920 0.525 3.620 ;
        RECT 3.605 2.920 3.835 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 4.910 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.605 0.300 3.835 0.930 ;
        RECT 0.000 -0.300 4.480 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.755 3.160 3.075 3.390 ;
        RECT 0.755 2.690 0.985 3.160 ;
        RECT 0.245 2.460 0.985 2.690 ;
        RECT 0.245 0.550 0.475 2.460 ;
        RECT 2.845 2.360 3.075 3.160 ;
        RECT 2.485 2.130 3.075 2.360 ;
        RECT 2.485 0.550 2.715 2.130 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai21_1
MACRO gf180mcu_fd_sc_mcu7t5v0__oai21_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai21_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.400 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.970 1.790 6.080 2.120 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.395 2.350 6.615 2.680 ;
        RECT 3.395 2.090 3.655 2.350 ;
        RECT 2.980 1.830 3.655 2.090 ;
        RECT 6.355 2.195 6.615 2.350 ;
        RECT 6.355 1.790 7.250 2.195 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.939000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.280 1.785 2.750 2.120 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.309600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 2.680 1.595 3.335 ;
        RECT 2.865 3.050 7.075 3.280 ;
        RECT 2.865 2.680 3.095 3.050 ;
        RECT 1.365 2.450 3.095 2.680 ;
        RECT 6.845 2.675 7.075 3.050 ;
        RECT 6.845 2.445 7.730 2.675 ;
        RECT 7.500 1.560 7.730 2.445 ;
        RECT 3.770 1.220 7.730 1.560 ;
        RECT 3.770 0.990 4.110 1.220 ;
        RECT 6.010 0.990 6.350 1.220 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 8.400 4.220 ;
        RECT 0.345 2.995 0.575 3.620 ;
        RECT 2.385 2.995 2.615 3.620 ;
        RECT 7.305 2.995 7.535 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 8.830 4.350 ;
        RECT -0.430 1.760 3.265 1.885 ;
        RECT 6.805 1.760 8.830 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.830 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 1.015 ;
        RECT 0.000 -0.300 8.400 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.310 2.715 1.545 ;
        RECT 0.245 0.635 0.475 1.310 ;
        RECT 2.485 0.760 2.715 1.310 ;
        RECT 2.485 0.530 7.700 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai21_2
MACRO gf180mcu_fd_sc_mcu7t5v0__oai21_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai21_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.120 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.530 1.800 3.580 2.120 ;
        RECT 3.350 1.680 3.580 1.800 ;
        RECT 3.350 1.450 8.070 1.680 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.680 2.360 4.100 2.680 ;
        RECT 0.680 1.695 1.000 2.360 ;
        RECT 3.870 2.140 4.100 2.360 ;
        RECT 3.870 1.910 9.140 2.140 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.878000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.020 1.800 14.550 2.120 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.030500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.085 3.055 4.640 3.240 ;
        RECT 5.480 3.055 9.615 3.240 ;
        RECT 1.085 2.920 9.615 3.055 ;
        RECT 4.410 2.825 5.710 2.920 ;
        RECT 9.385 2.680 9.615 2.920 ;
        RECT 10.865 2.680 11.095 3.250 ;
        RECT 12.905 2.680 13.135 3.250 ;
        RECT 9.385 2.360 13.135 2.680 ;
        RECT 9.385 1.220 9.615 2.360 ;
        RECT 1.520 0.990 9.615 1.220 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 15.120 4.220 ;
        RECT 0.245 2.910 0.475 3.620 ;
        RECT 4.890 3.285 5.230 3.620 ;
        RECT 9.845 2.910 10.075 3.620 ;
        RECT 11.885 2.910 12.115 3.620 ;
        RECT 13.925 2.910 14.155 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 15.550 4.350 ;
        RECT -0.430 1.760 1.140 1.885 ;
        RECT 10.055 1.760 15.550 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 15.550 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 10.765 0.300 10.995 0.910 ;
        RECT 13.005 0.300 13.235 0.910 ;
        RECT 0.000 -0.300 15.120 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 10.150 1.160 14.355 1.390 ;
        RECT 10.150 0.760 10.380 1.160 ;
        RECT 0.180 0.530 10.380 0.760 ;
        RECT 11.885 0.570 12.115 1.160 ;
        RECT 14.125 0.570 14.355 1.160 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai21_4
MACRO gf180mcu_fd_sc_mcu7t5v0__oai22_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai22_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.945 0.550 3.240 2.220 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.065 0.550 4.380 2.220 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 2.190 2.160 2.845 ;
        RECT 1.800 1.685 2.715 2.190 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 1.610 1.030 3.320 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal1 ;
        RECT 2.440 2.680 3.835 2.910 ;
        RECT 3.480 0.550 3.835 2.680 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.600 4.220 ;
        RECT 0.245 2.590 0.475 3.620 ;
        RECT 4.625 2.960 4.855 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 6.030 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.635 ;
        RECT 0.000 -0.300 5.600 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.320 3.140 4.365 3.370 ;
        RECT 1.320 1.095 1.550 3.140 ;
        RECT 4.135 2.680 4.365 3.140 ;
        RECT 4.135 2.450 4.955 2.680 ;
        RECT 0.245 0.865 2.715 1.095 ;
        RECT 0.245 0.550 0.475 0.865 ;
        RECT 2.485 0.550 2.715 0.865 ;
        RECT 4.725 0.550 4.955 2.450 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai22_1
MACRO gf180mcu_fd_sc_mcu7t5v0__oai22_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai22_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.640 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.250 1.800 8.715 2.120 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.690 2.360 9.295 2.680 ;
        RECT 5.690 2.120 6.020 2.360 ;
        RECT 5.270 1.800 6.020 2.120 ;
        RECT 8.955 1.585 9.295 2.360 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.475 1.785 3.270 2.120 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.825 2.360 3.820 2.680 ;
        RECT 0.825 1.585 1.165 2.360 ;
        RECT 3.500 2.125 3.820 2.360 ;
        RECT 3.500 1.770 4.480 2.125 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.377400 ;
    PORT
      LAYER Metal1 ;
        RECT 2.175 2.920 4.385 3.240 ;
        RECT 4.110 2.680 4.385 2.920 ;
        RECT 5.195 2.920 7.865 3.240 ;
        RECT 5.195 2.680 5.445 2.920 ;
        RECT 4.110 2.360 5.445 2.680 ;
        RECT 4.755 1.560 5.015 2.360 ;
        RECT 4.755 1.240 8.590 1.560 ;
        RECT 6.010 0.990 6.350 1.240 ;
        RECT 8.250 0.990 8.590 1.240 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 10.640 4.220 ;
        RECT 0.345 2.590 0.575 3.620 ;
        RECT 4.725 2.975 4.955 3.620 ;
        RECT 9.545 2.590 9.775 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 11.070 4.350 ;
        RECT -0.430 1.760 5.605 1.885 ;
        RECT 8.985 1.760 11.070 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 11.070 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 0.815 ;
        RECT 3.605 0.300 3.835 0.815 ;
        RECT 0.000 -0.300 10.640 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 1.045 4.455 1.275 ;
        RECT 0.190 0.530 0.530 1.045 ;
        RECT 2.430 0.530 2.770 1.045 ;
        RECT 4.225 0.760 4.455 1.045 ;
        RECT 4.225 0.530 9.940 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai22_2
MACRO gf180mcu_fd_sc_mcu7t5v0__oai22_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai22_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.600 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.730 1.785 12.540 2.120 ;
        RECT 12.290 1.680 12.540 1.785 ;
        RECT 12.290 1.450 17.120 1.680 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.200 2.360 13.125 2.680 ;
        RECT 10.200 2.120 10.500 2.360 ;
        RECT 9.610 1.800 10.500 2.120 ;
        RECT 12.875 2.140 13.125 2.360 ;
        RECT 12.875 1.910 18.460 2.140 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.530 1.785 3.360 2.120 ;
        RECT 3.110 1.635 3.360 1.785 ;
        RECT 3.110 1.405 7.940 1.635 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.825 2.360 3.940 2.680 ;
        RECT 0.825 1.585 1.145 2.360 ;
        RECT 3.690 2.095 3.940 2.360 ;
        RECT 3.690 1.865 8.850 2.095 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.369000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.730 3.025 4.420 3.240 ;
        RECT 5.255 3.025 8.905 3.380 ;
        RECT 9.740 3.025 13.605 3.240 ;
        RECT 14.440 3.025 16.375 3.380 ;
        RECT 1.730 2.920 16.375 3.025 ;
        RECT 4.170 2.795 9.990 2.920 ;
        RECT 13.355 2.795 14.690 2.920 ;
        RECT 6.910 2.570 7.250 2.795 ;
        RECT 9.080 1.220 9.380 2.795 ;
        RECT 16.145 2.485 16.375 2.920 ;
        RECT 9.080 0.990 17.560 1.220 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 19.600 4.220 ;
        RECT 0.345 2.590 0.575 3.620 ;
        RECT 4.670 3.255 5.010 3.620 ;
        RECT 9.150 3.255 9.490 3.620 ;
        RECT 13.850 3.255 14.190 3.620 ;
        RECT 18.505 2.590 18.735 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 20.030 4.350 ;
        RECT -0.430 1.760 10.090 1.885 ;
        RECT 17.950 1.760 20.030 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 20.030 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.715 ;
        RECT 3.550 0.300 3.890 0.715 ;
        RECT 5.790 0.300 6.130 0.715 ;
        RECT 8.030 0.300 8.370 0.715 ;
        RECT 0.000 -0.300 19.600 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.190 0.945 8.840 1.175 ;
        RECT 0.190 0.550 0.530 0.945 ;
        RECT 2.430 0.550 2.770 0.945 ;
        RECT 4.670 0.550 5.010 0.945 ;
        RECT 6.910 0.550 7.250 0.945 ;
        RECT 8.610 0.760 8.840 0.945 ;
        RECT 8.610 0.530 18.900 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai22_4
MACRO gf180mcu_fd_sc_mcu7t5v0__oai31_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai31_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.160 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.036500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.230 1.750 2.130 2.150 ;
        RECT 1.790 1.160 2.130 1.750 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.036500 ;
    PORT
      LAYER Metal1 ;
        RECT 3.470 1.470 3.810 3.320 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.036500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.590 1.470 4.935 3.320 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.054000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 1.160 1.000 3.320 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.988400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.330 2.680 1.670 3.380 ;
        RECT 1.330 2.380 2.680 2.680 ;
        RECT 2.360 1.220 2.680 2.380 ;
        RECT 2.360 0.990 5.395 1.220 ;
        RECT 5.165 0.605 5.395 0.990 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 6.160 4.220 ;
        RECT 0.245 2.530 0.475 3.620 ;
        RECT 5.165 2.530 5.395 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 6.590 4.350 ;
        RECT -0.430 1.760 2.195 1.885 ;
        RECT 3.440 1.760 6.590 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.590 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 0.945 ;
        RECT 0.000 -0.300 6.160 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.310 0.530 4.330 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai31_1
MACRO gf180mcu_fd_sc_mcu7t5v0__oai31_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai31_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.640 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.420 1.680 6.975 1.985 ;
        RECT 9.620 1.680 9.980 2.280 ;
        RECT 5.420 1.665 9.980 1.680 ;
        RECT 6.745 1.450 9.980 1.665 ;
        RECT 8.970 1.210 9.980 1.450 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 7.255 2.465 8.350 2.690 ;
        RECT 4.460 2.235 8.350 2.465 ;
        RECT 4.460 2.150 4.990 2.235 ;
        RECT 4.030 1.770 4.990 2.150 ;
        RECT 7.670 1.910 8.350 2.235 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.600 2.930 9.240 3.260 ;
        RECT 3.470 2.920 9.240 2.930 ;
        RECT 3.470 2.695 6.850 2.920 ;
        RECT 3.470 2.120 3.800 2.695 ;
        RECT 2.970 1.770 3.800 2.120 ;
        RECT 9.010 1.910 9.240 2.920 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.064000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.280 1.770 2.130 2.150 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.796000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 2.760 1.595 3.375 ;
        RECT 2.970 3.160 6.350 3.390 ;
        RECT 2.970 2.760 3.200 3.160 ;
        RECT 1.365 2.530 3.200 2.760 ;
        RECT 2.360 1.220 2.680 2.530 ;
        RECT 2.360 0.990 8.600 1.220 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 10.640 4.220 ;
        RECT 0.295 2.530 0.525 3.620 ;
        RECT 2.330 3.020 2.670 3.620 ;
        RECT 9.490 2.530 9.830 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 11.070 4.350 ;
        RECT -0.430 1.760 3.340 1.885 ;
        RECT 9.070 1.760 11.070 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 11.070 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.635 ;
        RECT 0.000 -0.300 10.640 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.180 0.865 2.130 1.095 ;
        RECT 1.900 0.760 2.130 0.865 ;
        RECT 1.900 0.530 9.940 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai31_2
MACRO gf180mcu_fd_sc_mcu7t5v0__oai31_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai31_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.600 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.480 1.770 4.920 2.150 ;
        RECT 4.690 1.680 4.920 1.770 ;
        RECT 4.690 1.450 12.420 1.680 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.150 2.450 6.775 2.710 ;
        RECT 5.150 2.220 13.890 2.450 ;
        RECT 5.420 1.910 5.920 2.220 ;
        RECT 8.860 1.910 10.220 2.220 ;
        RECT 12.970 1.725 13.890 2.220 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.620 1.680 3.240 2.150 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.890 1.785 19.150 2.120 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.028900 ;
    PORT
      LAYER Metal1 ;
        RECT 7.130 2.700 18.430 2.930 ;
        RECT 14.120 2.360 18.430 2.700 ;
        RECT 14.120 1.220 14.440 2.360 ;
        RECT 1.310 0.990 14.440 1.220 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 19.600 4.220 ;
        RECT 1.530 3.285 1.870 3.620 ;
        RECT 3.770 3.285 4.110 3.620 ;
        RECT 14.470 3.285 14.810 3.620 ;
        RECT 16.610 3.285 16.950 3.620 ;
        RECT 18.855 2.570 19.085 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 20.030 4.350 ;
        RECT -0.430 1.760 1.095 1.885 ;
        RECT 14.580 1.760 20.030 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 20.030 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 15.490 0.300 15.830 0.635 ;
        RECT 17.730 0.300 18.070 0.635 ;
        RECT 0.000 -0.300 19.600 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 2.800 0.575 3.380 ;
        RECT 2.705 2.800 2.935 3.380 ;
        RECT 4.360 3.160 14.100 3.390 ;
        RECT 4.360 2.800 4.590 3.160 ;
        RECT 0.345 2.570 4.590 2.800 ;
        RECT 14.980 0.865 19.200 1.095 ;
        RECT 14.980 0.760 15.210 0.865 ;
        RECT 0.180 0.530 15.210 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai31_4
MACRO gf180mcu_fd_sc_mcu7t5v0__oai32_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai32_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.920 2.150 3.240 2.750 ;
        RECT 2.920 1.730 3.830 2.150 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 1.650 2.120 3.310 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 1.650 1.000 3.310 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.065 0.610 4.370 2.150 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.185 0.610 5.490 2.190 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.304800 ;
    PORT
      LAYER Metal1 ;
        RECT 3.470 2.380 4.955 2.700 ;
        RECT 4.600 0.610 4.955 2.380 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 6.720 4.220 ;
        RECT 0.245 2.590 0.475 3.620 ;
        RECT 5.745 3.200 5.975 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 7.150 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.150 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 0.915 ;
        RECT 2.485 0.300 2.715 0.915 ;
        RECT 0.000 -0.300 6.720 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.450 3.050 5.450 3.280 ;
        RECT 2.450 1.400 2.680 3.050 ;
        RECT 5.220 2.870 5.450 3.050 ;
        RECT 5.220 2.640 6.075 2.870 ;
        RECT 1.365 1.165 3.835 1.400 ;
        RECT 1.365 0.610 1.595 1.165 ;
        RECT 3.605 0.610 3.835 1.165 ;
        RECT 5.845 0.610 6.075 2.640 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai32_1
MACRO gf180mcu_fd_sc_mcu7t5v0__oai32_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai32_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.880 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.850 1.800 4.390 2.120 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.535 1.770 2.600 2.135 ;
        RECT 2.350 1.555 2.600 1.770 ;
        RECT 4.620 1.770 6.070 2.120 ;
        RECT 4.620 1.555 4.850 1.770 ;
        RECT 2.350 1.325 4.850 1.555 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.825 2.595 6.160 2.680 ;
        RECT 0.825 2.365 6.600 2.595 ;
        RECT 0.825 1.560 1.145 2.365 ;
        RECT 6.300 1.560 6.600 2.365 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.450 1.800 10.590 2.120 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.120 2.595 11.535 2.680 ;
        RECT 7.560 2.365 11.535 2.595 ;
        RECT 7.560 1.785 7.880 2.365 ;
        RECT 11.215 1.560 11.535 2.365 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.377400 ;
    PORT
      LAYER Metal1 ;
        RECT 3.365 3.055 6.660 3.240 ;
        RECT 7.500 3.055 10.170 3.240 ;
        RECT 3.365 2.920 10.170 3.055 ;
        RECT 6.410 2.825 7.750 2.920 ;
        RECT 6.840 1.220 7.160 2.825 ;
        RECT 6.840 0.990 10.840 1.220 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 12.880 4.220 ;
        RECT 0.345 2.650 0.575 3.620 ;
        RECT 6.910 3.285 7.250 3.620 ;
        RECT 11.785 2.650 12.015 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 13.310 4.350 ;
        RECT -0.430 1.760 7.770 1.885 ;
        RECT 11.280 1.760 13.310 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.310 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.635 ;
        RECT 3.550 0.300 3.890 0.635 ;
        RECT 5.790 0.300 6.130 0.635 ;
        RECT 0.000 -0.300 12.880 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.180 0.865 6.600 1.095 ;
        RECT 6.370 0.760 6.600 0.865 ;
        RECT 6.370 0.530 12.180 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai32_2
MACRO gf180mcu_fd_sc_mcu7t5v0__oai32_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai32_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.080 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.570 1.800 13.880 2.120 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.730 2.580 6.365 2.690 ;
        RECT 1.055 2.350 9.135 2.580 ;
        RECT 1.055 1.760 1.295 2.350 ;
        RECT 4.365 1.825 5.725 2.350 ;
        RECT 8.895 1.760 9.135 2.350 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.730 1.800 3.870 2.120 ;
        RECT 3.640 1.575 3.870 1.800 ;
        RECT 6.210 1.800 8.350 2.120 ;
        RECT 6.210 1.575 6.440 1.800 ;
        RECT 3.640 1.345 6.440 1.575 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 16.005 1.800 17.870 2.120 ;
        RECT 17.640 1.680 17.870 1.800 ;
        RECT 20.210 1.800 22.350 2.120 ;
        RECT 20.210 1.680 20.440 1.800 ;
        RECT 17.640 1.450 20.440 1.680 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.545 2.595 18.050 2.680 ;
        RECT 19.945 2.595 23.225 2.680 ;
        RECT 15.545 2.360 23.225 2.595 ;
        RECT 15.545 2.120 15.775 2.360 ;
        RECT 14.650 1.800 15.775 2.120 ;
        RECT 18.325 1.910 19.685 2.360 ;
        RECT 22.965 1.760 23.225 2.360 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.176100 ;
    PORT
      LAYER Metal1 ;
        RECT 15.045 3.055 18.585 3.240 ;
        RECT 19.425 3.055 21.810 3.240 ;
        RECT 15.045 2.920 21.810 3.055 ;
        RECT 15.045 2.815 15.295 2.920 ;
        RECT 18.335 2.825 19.655 2.920 ;
        RECT 9.570 2.360 15.295 2.815 ;
        RECT 14.120 1.220 14.420 2.360 ;
        RECT 14.120 0.990 22.535 1.220 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 24.080 4.220 ;
        RECT 2.635 3.285 2.975 3.620 ;
        RECT 7.115 3.285 7.455 3.620 ;
        RECT 14.455 3.285 14.795 3.620 ;
        RECT 18.835 3.285 19.175 3.620 ;
        RECT 23.500 2.530 23.730 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 24.510 4.350 ;
        RECT -0.430 1.760 13.825 1.885 ;
        RECT 22.980 1.760 24.510 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 24.510 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.515 0.300 1.855 0.635 ;
        RECT 3.755 0.300 4.095 0.635 ;
        RECT 5.995 0.300 6.335 0.635 ;
        RECT 8.235 0.300 8.575 0.635 ;
        RECT 10.475 0.300 10.815 0.635 ;
        RECT 12.715 0.300 13.055 0.635 ;
        RECT 0.000 -0.300 24.080 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.500 3.055 0.730 3.380 ;
        RECT 3.230 3.055 6.865 3.170 ;
        RECT 8.190 3.140 14.085 3.370 ;
        RECT 8.190 3.055 8.420 3.140 ;
        RECT 0.500 2.940 8.420 3.055 ;
        RECT 0.500 2.825 3.480 2.940 ;
        RECT 6.615 2.825 8.420 2.940 ;
        RECT 0.500 2.530 0.730 2.825 ;
        RECT 0.385 0.865 13.635 1.095 ;
        RECT 13.405 0.760 13.635 0.865 ;
        RECT 13.405 0.530 23.885 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai32_4
MACRO gf180mcu_fd_sc_mcu7t5v0__oai33_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai33_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.400 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.039500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.040 1.525 4.360 3.320 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.039500 ;
    PORT
      LAYER Metal1 ;
        RECT 5.160 2.140 5.480 3.320 ;
        RECT 5.160 1.770 6.040 2.140 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.039500 ;
    PORT
      LAYER Metal1 ;
        RECT 6.280 2.140 6.600 3.320 ;
        RECT 6.280 1.770 7.870 2.140 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.039500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.920 1.525 3.240 3.320 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.039500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 1.525 2.120 3.320 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.039500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 1.525 1.000 3.320 ;
    END
  END B3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.871900 ;
    PORT
      LAYER Metal1 ;
        RECT 3.490 1.220 3.790 3.380 ;
        RECT 3.490 0.990 7.635 1.220 ;
        RECT 7.405 0.555 7.635 0.990 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 8.400 4.220 ;
        RECT 0.245 2.530 0.475 3.620 ;
        RECT 7.305 2.530 7.535 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 8.830 4.350 ;
        RECT -0.430 1.760 4.410 1.885 ;
        RECT 5.695 1.760 8.830 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.830 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 0.815 ;
        RECT 2.485 0.300 2.715 0.815 ;
        RECT 0.000 -0.300 8.400 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 1.045 3.175 1.275 ;
        RECT 1.365 0.530 1.595 1.045 ;
        RECT 2.945 0.760 3.175 1.045 ;
        RECT 2.945 0.530 6.570 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai33_1
MACRO gf180mcu_fd_sc_mcu7t5v0__oai33_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai33_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.120 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.120 1.680 14.440 2.380 ;
        RECT 9.800 1.450 14.440 1.680 ;
        RECT 13.380 1.160 14.440 1.450 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.480 1.910 12.540 2.140 ;
        RECT 8.480 1.780 9.520 1.910 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.000 2.370 13.775 2.680 ;
        RECT 8.000 2.140 8.230 2.370 ;
        RECT 7.440 1.780 8.230 2.140 ;
        RECT 13.435 1.910 13.775 2.370 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.890 1.800 4.950 2.120 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.510 1.770 2.660 2.150 ;
        RECT 2.410 1.555 2.660 1.770 ;
        RECT 5.180 1.555 5.480 2.150 ;
        RECT 2.410 1.325 5.480 1.555 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.825 2.380 6.060 2.680 ;
        RECT 0.825 2.120 1.145 2.380 ;
        RECT 0.280 1.800 1.145 2.120 ;
        RECT 5.720 2.120 6.060 2.380 ;
        RECT 5.720 1.800 6.600 2.120 ;
    END
  END B3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.803800 ;
    PORT
      LAYER Metal1 ;
        RECT 2.750 3.055 6.660 3.240 ;
        RECT 7.500 3.055 11.215 3.240 ;
        RECT 2.750 2.920 11.215 3.055 ;
        RECT 6.410 2.825 7.750 2.920 ;
        RECT 6.850 1.220 7.150 2.825 ;
        RECT 6.850 0.990 13.070 1.220 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 15.120 4.220 ;
        RECT 0.345 2.630 0.575 3.620 ;
        RECT 6.910 3.285 7.250 3.620 ;
        RECT 14.025 2.630 14.255 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 15.550 4.350 ;
        RECT -0.430 1.760 7.800 1.885 ;
        RECT 13.565 1.760 15.550 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 15.550 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.635 ;
        RECT 3.550 0.300 3.890 0.635 ;
        RECT 5.790 0.300 6.130 0.635 ;
        RECT 0.000 -0.300 15.120 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.180 0.865 6.610 1.095 ;
        RECT 6.380 0.760 6.610 0.865 ;
        RECT 6.380 0.530 14.420 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai33_2
MACRO gf180mcu_fd_sc_mcu7t5v0__oai33_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai33_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.560 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 14.580 1.800 18.440 2.120 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 21.955 2.590 24.605 2.710 ;
        RECT 19.290 2.360 27.490 2.590 ;
        RECT 19.290 1.760 19.530 2.360 ;
        RECT 22.600 1.920 23.960 2.360 ;
        RECT 27.250 1.760 27.490 2.360 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 20.180 1.800 21.915 2.120 ;
        RECT 21.685 1.680 21.915 1.800 ;
        RECT 24.545 1.800 26.835 2.120 ;
        RECT 24.545 1.680 24.775 1.800 ;
        RECT 21.685 1.450 24.775 1.680 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.580 1.800 13.340 2.120 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.520 2.595 6.160 2.700 ;
        RECT 0.775 2.360 8.840 2.595 ;
        RECT 0.775 1.530 1.095 2.360 ;
        RECT 4.160 1.920 5.520 2.360 ;
        RECT 8.580 1.760 8.840 2.360 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.740 1.800 3.820 2.120 ;
        RECT 3.590 1.565 3.820 1.800 ;
        RECT 6.220 1.800 8.310 2.120 ;
        RECT 6.220 1.565 6.450 1.800 ;
        RECT 3.590 1.335 6.450 1.565 ;
    END
  END B3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.028900 ;
    PORT
      LAYER Metal1 ;
        RECT 9.580 2.360 17.890 2.795 ;
        RECT 13.570 1.220 13.870 2.360 ;
        RECT 13.570 0.990 26.820 1.220 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 28.560 4.220 ;
        RECT 2.430 3.285 2.770 3.620 ;
        RECT 6.910 3.285 7.250 3.620 ;
        RECT 20.870 3.285 21.210 3.620 ;
        RECT 25.350 3.285 25.690 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 28.990 4.350 ;
        RECT -0.430 1.760 13.550 1.885 ;
        RECT 27.235 1.760 28.990 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 28.990 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.635 ;
        RECT 3.550 0.300 3.890 0.635 ;
        RECT 5.790 0.300 6.130 0.635 ;
        RECT 8.030 0.300 8.370 0.635 ;
        RECT 10.270 0.300 10.610 0.635 ;
        RECT 12.510 0.300 12.850 0.635 ;
        RECT 0.000 -0.300 28.560 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.295 3.055 0.525 3.380 ;
        RECT 3.020 3.090 6.660 3.320 ;
        RECT 3.020 3.055 3.270 3.090 ;
        RECT 0.295 2.825 3.270 3.055 ;
        RECT 6.410 3.055 6.660 3.090 ;
        RECT 7.500 3.090 13.870 3.320 ;
        RECT 14.240 3.090 20.355 3.320 ;
        RECT 7.500 3.055 7.730 3.090 ;
        RECT 6.410 2.825 7.730 3.055 ;
        RECT 20.110 3.055 20.355 3.090 ;
        RECT 21.460 3.090 25.100 3.320 ;
        RECT 21.460 3.055 21.705 3.090 ;
        RECT 20.110 2.825 21.705 3.055 ;
        RECT 24.855 3.055 25.100 3.090 ;
        RECT 27.765 3.055 27.995 3.380 ;
        RECT 24.855 2.825 27.995 3.055 ;
        RECT 0.295 2.530 0.525 2.825 ;
        RECT 27.765 2.530 27.995 2.825 ;
        RECT 0.180 0.865 13.330 1.095 ;
        RECT 13.100 0.760 13.330 0.865 ;
        RECT 13.100 0.530 28.160 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai33_4
MACRO gf180mcu_fd_sc_mcu7t5v0__oai211_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai211_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.825 0.550 2.120 2.135 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 0.550 1.000 2.230 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.984500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.360 1.800 3.370 2.120 ;
        RECT 2.360 1.160 2.660 1.800 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.984500 ;
    PORT
      LAYER Metal1 ;
        RECT 3.650 1.800 4.970 2.120 ;
        RECT 3.650 1.560 3.940 1.800 ;
        RECT 2.890 1.240 3.940 1.560 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.672850 ;
    PORT
      LAYER Metal1 ;
        RECT 2.430 2.700 2.770 2.930 ;
        RECT 1.240 2.595 2.770 2.700 ;
        RECT 4.580 2.595 4.920 2.930 ;
        RECT 1.240 2.365 4.920 2.595 ;
        RECT 1.240 0.550 1.595 2.365 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.600 4.220 ;
        RECT 0.295 2.920 0.525 3.620 ;
        RECT 3.550 3.285 3.890 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 6.030 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 4.725 0.300 4.955 0.890 ;
        RECT 0.000 -0.300 5.600 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.755 3.160 3.290 3.390 ;
        RECT 0.755 2.690 0.985 3.160 ;
        RECT 3.060 3.055 3.290 3.160 ;
        RECT 4.120 3.160 5.450 3.390 ;
        RECT 4.120 3.055 4.350 3.160 ;
        RECT 3.060 2.825 4.350 3.055 ;
        RECT 0.245 2.460 0.985 2.690 ;
        RECT 0.245 0.550 0.475 2.460 ;
        RECT 5.220 1.370 5.450 3.160 ;
        RECT 4.240 1.140 5.450 1.370 ;
        RECT 4.240 0.835 4.470 1.140 ;
        RECT 2.430 0.605 4.470 0.835 ;
        RECT 4.240 0.600 4.470 0.605 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai211_1
MACRO gf180mcu_fd_sc_mcu7t5v0__oai211_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai211_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.560 1.790 3.870 2.120 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.825 2.350 4.380 2.680 ;
        RECT 0.825 1.160 1.145 2.350 ;
        RECT 4.120 2.120 4.380 2.350 ;
        RECT 4.120 1.790 4.900 2.120 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.969000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.720 1.555 6.040 2.150 ;
        RECT 8.865 1.555 9.420 2.190 ;
        RECT 5.720 1.325 9.420 1.555 ;
        RECT 5.720 1.190 6.485 1.325 ;
        RECT 8.380 1.190 9.420 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.969000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.280 1.800 8.320 2.140 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.837400 ;
    PORT
      LAYER Metal1 ;
        RECT 2.130 2.920 4.860 3.280 ;
        RECT 4.630 2.680 4.860 2.920 ;
        RECT 6.290 2.680 6.520 3.275 ;
        RECT 8.330 2.680 8.560 3.275 ;
        RECT 4.630 2.380 8.560 2.680 ;
        RECT 4.630 2.370 5.480 2.380 ;
        RECT 5.150 1.560 5.480 2.370 ;
        RECT 1.530 1.220 5.480 1.560 ;
        RECT 1.530 0.990 1.870 1.220 ;
        RECT 3.770 0.990 4.110 1.220 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 10.080 4.220 ;
        RECT 0.345 2.485 0.575 3.620 ;
        RECT 5.115 3.205 5.455 3.620 ;
        RECT 7.255 3.205 7.595 3.620 ;
        RECT 9.350 2.595 9.580 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 10.510 4.350 ;
        RECT -0.430 1.760 1.075 1.885 ;
        RECT 4.615 1.760 10.510 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 7.255 0.300 7.595 0.635 ;
        RECT 0.000 -0.300 10.080 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 6.735 0.865 8.080 1.095 ;
        RECT 6.735 0.760 6.965 0.865 ;
        RECT 0.180 0.530 6.965 0.760 ;
        RECT 7.850 0.760 8.080 0.865 ;
        RECT 7.850 0.530 9.645 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai211_2
MACRO gf180mcu_fd_sc_mcu7t5v0__oai211_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai211_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.480 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.540 1.770 8.310 2.120 ;
        RECT 6.540 1.680 6.790 1.770 ;
        RECT 1.960 1.450 6.790 1.680 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.955 2.360 8.880 2.680 ;
        RECT 5.955 2.140 6.205 2.360 ;
        RECT 0.620 1.910 6.205 2.140 ;
        RECT 8.540 2.120 8.880 2.360 ;
        RECT 8.540 1.770 9.410 2.120 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.938000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.200 1.555 10.520 2.425 ;
        RECT 10.200 1.325 17.760 1.555 ;
        RECT 12.930 1.220 15.080 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.938000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.750 1.800 16.840 2.120 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.279000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.650 3.240 2.990 3.325 ;
        RECT 2.650 3.025 4.640 3.240 ;
        RECT 5.475 3.025 9.340 3.240 ;
        RECT 10.175 3.055 11.480 3.240 ;
        RECT 12.320 3.055 13.520 3.240 ;
        RECT 14.360 3.055 15.560 3.240 ;
        RECT 16.400 3.055 17.450 3.240 ;
        RECT 10.175 3.025 17.450 3.055 ;
        RECT 2.650 2.920 17.450 3.025 ;
        RECT 2.650 2.475 2.990 2.920 ;
        RECT 4.390 2.795 5.725 2.920 ;
        RECT 9.090 2.795 17.450 2.920 ;
        RECT 9.640 1.220 9.960 2.795 ;
        RECT 1.520 0.990 9.960 1.220 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 18.480 4.220 ;
        RECT 0.345 2.530 0.575 3.620 ;
        RECT 4.890 3.285 5.230 3.620 ;
        RECT 9.590 3.285 9.930 3.620 ;
        RECT 11.730 3.285 12.070 3.620 ;
        RECT 13.770 3.285 14.110 3.620 ;
        RECT 15.810 3.285 16.150 3.620 ;
        RECT 17.905 2.595 18.135 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 18.910 4.350 ;
        RECT -0.430 1.760 1.135 1.885 ;
        RECT 8.995 1.760 18.910 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.910 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 11.730 0.300 12.070 0.635 ;
        RECT 15.810 0.300 16.150 0.635 ;
        RECT 0.000 -0.300 18.480 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 10.655 0.865 12.550 1.095 ;
        RECT 10.655 0.760 10.885 0.865 ;
        RECT 0.180 0.530 10.885 0.760 ;
        RECT 12.320 0.760 12.550 0.865 ;
        RECT 15.330 0.865 18.200 1.095 ;
        RECT 15.330 0.760 15.560 0.865 ;
        RECT 12.320 0.530 15.560 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai211_4
MACRO gf180mcu_fd_sc_mcu7t5v0__oai221_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai221_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.160 1.770 6.110 2.150 ;
        RECT 5.160 1.170 5.500 1.770 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.010 1.170 4.390 2.135 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.240 1.575 1.560 3.320 ;
        RECT 1.240 1.345 2.110 1.575 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 1.345 1.000 3.320 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.964500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.340 1.210 3.260 1.665 ;
        RECT 2.945 0.610 3.260 1.210 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.753600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.430 2.595 2.770 2.930 ;
        RECT 5.770 2.700 6.110 2.930 ;
        RECT 4.795 2.595 6.110 2.700 ;
        RECT 2.430 2.380 6.110 2.595 ;
        RECT 2.430 2.365 4.910 2.380 ;
        RECT 4.620 0.910 4.910 2.365 ;
        RECT 4.620 0.610 5.095 0.910 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 6.720 4.220 ;
        RECT 0.245 2.530 0.475 3.620 ;
        RECT 3.610 3.285 3.950 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 7.150 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.150 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.635 ;
        RECT 0.000 -0.300 6.720 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.950 3.160 3.360 3.390 ;
        RECT 1.950 2.135 2.180 3.160 ;
        RECT 3.130 3.055 3.360 3.160 ;
        RECT 4.290 3.160 6.570 3.390 ;
        RECT 4.290 3.055 4.520 3.160 ;
        RECT 3.130 2.825 4.520 3.055 ;
        RECT 1.950 1.905 3.770 2.135 ;
        RECT 0.245 0.965 2.110 1.095 ;
        RECT 0.245 0.865 2.715 0.965 ;
        RECT 0.245 0.625 0.475 0.865 ;
        RECT 1.880 0.625 2.715 0.865 ;
        RECT 3.540 0.910 3.770 1.905 ;
        RECT 6.340 0.910 6.570 3.160 ;
        RECT 3.540 0.680 3.950 0.910 ;
        RECT 5.870 0.680 6.570 0.910 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai221_1
MACRO gf180mcu_fd_sc_mcu7t5v0__oai221_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai221_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.880 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.550 2.365 11.570 2.595 ;
        RECT 8.550 2.150 8.820 2.365 ;
        RECT 8.160 1.770 8.820 2.150 ;
        RECT 11.340 2.150 11.570 2.365 ;
        RECT 11.340 1.770 12.590 2.150 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 9.050 1.800 11.110 2.120 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.530 1.800 4.710 2.120 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.625 1.570 1.000 2.275 ;
        RECT 0.625 1.340 4.455 1.570 ;
        RECT 0.625 1.160 1.690 1.340 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.969000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.105 1.800 7.330 2.120 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.382000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.485 2.680 2.715 3.375 ;
        RECT 5.545 2.680 5.775 3.110 ;
        RECT 7.560 3.055 9.540 3.260 ;
        RECT 10.525 3.055 12.580 3.260 ;
        RECT 7.560 2.825 12.580 3.055 ;
        RECT 7.560 2.680 7.915 2.825 ;
        RECT 2.485 2.360 7.915 2.680 ;
        RECT 7.560 1.220 7.915 2.360 ;
        RECT 7.560 0.990 11.330 1.220 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 12.880 4.220 ;
        RECT 0.245 2.690 0.475 3.620 ;
        RECT 4.670 3.090 5.010 3.620 ;
        RECT 6.510 3.090 6.850 3.620 ;
        RECT 9.870 3.285 10.210 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 13.310 4.350 ;
        RECT -0.430 1.760 4.965 1.885 ;
        RECT 11.780 1.760 13.310 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.310 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.185 0.300 0.530 0.635 ;
        RECT 2.425 0.300 2.770 0.635 ;
        RECT 4.665 0.300 5.010 0.635 ;
        RECT 0.000 -0.300 12.880 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 4.860 1.095 6.865 1.220 ;
        RECT 1.940 0.990 6.865 1.095 ;
        RECT 1.940 0.865 5.110 0.990 ;
        RECT 1.940 0.780 2.170 0.865 ;
        RECT 1.260 0.550 2.170 0.780 ;
        RECT 5.380 0.530 12.680 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai221_2
MACRO gf180mcu_fd_sc_mcu7t5v0__oai221_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai221_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.080 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 17.970 2.595 20.110 2.680 ;
        RECT 15.015 2.365 20.110 2.595 ;
        RECT 15.015 1.600 15.245 2.365 ;
        RECT 18.320 1.910 18.660 2.365 ;
        RECT 19.340 2.140 20.110 2.365 ;
        RECT 19.340 1.910 23.420 2.140 ;
        RECT 22.385 1.790 23.420 1.910 ;
        RECT 23.060 1.120 23.420 1.790 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.715 1.800 17.925 2.120 ;
        RECT 17.675 1.680 17.925 1.800 ;
        RECT 17.675 1.450 21.880 1.680 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.620 1.800 1.590 2.120 ;
        RECT 1.350 1.570 1.590 1.800 ;
        RECT 7.940 1.770 9.470 2.120 ;
        RECT 7.940 1.570 8.170 1.770 ;
        RECT 1.350 1.340 8.170 1.570 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.840 1.800 7.710 2.120 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.838000 ;
    PORT
      LAYER Metal1 ;
        RECT 10.115 1.800 14.160 2.120 ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.744200 ;
    PORT
      LAYER Metal1 ;
        RECT 0.345 2.680 0.575 3.110 ;
        RECT 4.725 2.680 4.955 3.110 ;
        RECT 9.205 2.680 9.435 3.110 ;
        RECT 10.025 2.680 10.255 3.110 ;
        RECT 12.165 2.680 12.395 3.110 ;
        RECT 17.235 3.055 20.735 3.310 ;
        RECT 14.350 2.910 23.780 3.055 ;
        RECT 14.350 2.825 17.465 2.910 ;
        RECT 20.505 2.825 23.780 2.910 ;
        RECT 14.350 2.680 14.690 2.825 ;
        RECT 0.345 2.360 14.690 2.680 ;
        RECT 14.405 1.220 14.690 2.360 ;
        RECT 14.405 0.990 22.530 1.220 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 24.080 4.220 ;
        RECT 2.430 3.090 2.770 3.620 ;
        RECT 6.910 3.090 7.250 3.620 ;
        RECT 10.990 3.090 11.330 3.620 ;
        RECT 13.230 3.090 13.570 3.620 ;
        RECT 16.590 3.285 16.930 3.620 ;
        RECT 21.070 3.285 21.410 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 24.510 4.350 ;
        RECT -0.430 1.760 9.445 1.885 ;
        RECT 22.940 1.760 24.510 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 24.510 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 0.635 ;
        RECT 2.425 0.300 2.770 0.635 ;
        RECT 4.665 0.300 5.010 0.635 ;
        RECT 6.905 0.300 7.250 0.635 ;
        RECT 9.145 0.300 9.490 0.635 ;
        RECT 0.000 -0.300 24.080 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 8.785 1.095 13.570 1.220 ;
        RECT 1.220 0.990 13.570 1.095 ;
        RECT 1.220 0.865 9.035 0.990 ;
        RECT 9.860 0.530 23.880 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai221_4
MACRO gf180mcu_fd_sc_mcu7t5v0__oai222_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai222_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.400 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.039500 ;
    PORT
      LAYER Metal1 ;
        RECT 7.300 1.770 8.270 2.150 ;
        RECT 7.300 1.060 7.720 1.770 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.039500 ;
    PORT
      LAYER Metal1 ;
        RECT 5.720 1.770 6.610 2.150 ;
        RECT 5.720 1.060 6.040 1.770 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.039500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.370 2.150 2.690 3.320 ;
        RECT 2.370 1.770 4.360 2.150 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.039500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.590 1.770 5.480 2.150 ;
        RECT 5.160 1.060 5.480 1.770 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.039500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.780 1.520 2.140 3.320 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.039500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.660 1.160 1.020 2.710 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.568400 ;
    PORT
      LAYER Metal1 ;
        RECT 3.055 2.970 5.065 3.260 ;
        RECT 6.035 2.970 8.100 3.260 ;
        RECT 3.055 2.900 8.100 2.970 ;
        RECT 4.755 2.740 8.100 2.900 ;
        RECT 6.840 1.220 7.070 2.740 ;
        RECT 6.510 0.990 7.070 1.220 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 8.400 4.220 ;
        RECT 0.345 2.950 0.575 3.620 ;
        RECT 5.445 3.200 5.675 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 8.830 4.350 ;
        RECT -0.430 1.760 2.725 1.885 ;
        RECT 7.300 1.760 8.830 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 2.725 1.760 7.300 1.885 ;
        RECT -0.430 -0.430 8.830 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 0.760 ;
        RECT 2.485 0.300 2.715 0.760 ;
        RECT 0.000 -0.300 8.400 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 0.990 4.610 1.220 ;
        RECT 1.365 0.530 1.595 0.990 ;
        RECT 3.150 0.530 8.200 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai222_1
MACRO gf180mcu_fd_sc_mcu7t5v0__oai222_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai222_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.120 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.285 2.595 14.460 2.690 ;
        RECT 10.525 2.365 14.460 2.595 ;
        RECT 10.525 1.645 11.060 2.365 ;
        RECT 14.005 1.160 14.460 2.365 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.290 1.800 13.390 2.120 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.070 2.595 6.740 2.690 ;
        RECT 5.070 2.365 9.380 2.595 ;
        RECT 6.040 1.790 6.300 2.365 ;
        RECT 9.100 2.150 9.380 2.365 ;
        RECT 9.100 1.770 9.680 2.150 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 6.770 1.800 8.870 2.120 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.660 1.570 1.020 2.190 ;
        RECT 4.010 1.800 5.015 2.120 ;
        RECT 4.010 1.570 4.380 1.800 ;
        RECT 0.660 1.335 4.380 1.570 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.530 1.800 3.460 2.120 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.265000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.125 3.055 7.340 3.240 ;
        RECT 8.445 3.055 11.775 3.240 ;
        RECT 12.720 3.055 14.820 3.240 ;
        RECT 0.280 2.920 14.820 3.055 ;
        RECT 0.280 2.825 3.420 2.920 ;
        RECT 7.090 2.825 12.950 2.920 ;
        RECT 9.930 1.220 10.160 2.825 ;
        RECT 9.930 0.990 13.570 1.220 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 15.120 4.220 ;
        RECT 2.430 3.285 2.770 3.620 ;
        RECT 7.630 3.285 7.970 3.620 ;
        RECT 12.110 3.285 12.450 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 15.550 4.350 ;
        RECT -0.430 1.760 4.940 1.885 ;
        RECT 13.995 1.760 15.550 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 15.550 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 0.845 ;
        RECT 2.430 0.300 2.770 0.635 ;
        RECT 4.670 0.300 5.010 0.635 ;
        RECT 0.000 -0.300 15.120 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 4.880 1.095 9.090 1.220 ;
        RECT 1.310 0.990 9.090 1.095 ;
        RECT 1.310 0.865 5.130 0.990 ;
        RECT 5.390 0.530 14.920 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai222_2
MACRO gf180mcu_fd_sc_mcu7t5v0__oai222_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai222_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.560 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 22.160 2.580 24.800 2.680 ;
        RECT 19.490 2.350 27.715 2.580 ;
        RECT 19.490 1.790 19.730 2.350 ;
        RECT 22.800 1.950 23.140 2.350 ;
        RECT 23.820 1.950 24.160 2.350 ;
        RECT 27.420 1.720 27.715 2.350 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 20.210 1.800 22.350 2.120 ;
        RECT 22.070 1.700 22.350 1.800 ;
        RECT 24.690 1.800 26.830 2.120 ;
        RECT 24.690 1.700 24.970 1.800 ;
        RECT 22.070 1.470 24.970 1.700 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.200 2.580 15.840 2.680 ;
        RECT 10.860 2.350 18.560 2.580 ;
        RECT 10.860 2.150 11.090 2.350 ;
        RECT 9.630 1.770 11.090 2.150 ;
        RECT 13.840 1.950 14.180 2.350 ;
        RECT 14.860 1.950 15.200 2.350 ;
        RECT 18.220 1.950 18.560 2.350 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 11.320 1.800 13.390 2.120 ;
        RECT 12.930 1.700 13.390 1.800 ;
        RECT 15.620 1.800 17.870 2.120 ;
        RECT 15.620 1.700 15.850 1.800 ;
        RECT 12.930 1.470 15.850 1.700 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.280 1.770 1.570 2.150 ;
        RECT 1.255 1.560 1.570 1.770 ;
        RECT 8.200 1.770 9.400 2.150 ;
        RECT 8.200 1.560 8.515 1.770 ;
        RECT 1.255 1.330 8.515 1.560 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.920 1.800 7.840 2.120 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.880750 ;
    PORT
      LAYER Metal1 ;
        RECT 0.295 3.050 0.525 3.380 ;
        RECT 4.725 3.240 4.955 3.380 ;
        RECT 3.020 3.050 6.660 3.240 ;
        RECT 12.700 3.050 16.340 3.240 ;
        RECT 18.810 3.050 19.120 3.380 ;
        RECT 21.660 3.050 25.300 3.240 ;
        RECT 27.965 3.050 28.195 3.380 ;
        RECT 0.295 2.920 28.195 3.050 ;
        RECT 0.295 2.820 12.950 2.920 ;
        RECT 16.090 2.820 21.910 2.920 ;
        RECT 25.050 2.820 28.195 2.920 ;
        RECT 0.295 2.530 0.525 2.820 ;
        RECT 4.725 2.530 4.955 2.820 ;
        RECT 18.810 1.220 19.120 2.820 ;
        RECT 27.965 2.530 28.195 2.820 ;
        RECT 18.810 0.990 27.010 1.220 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 28.560 4.220 ;
        RECT 2.430 3.280 2.770 3.620 ;
        RECT 6.910 3.285 7.250 3.620 ;
        RECT 12.110 3.285 12.450 3.620 ;
        RECT 16.590 3.285 16.930 3.620 ;
        RECT 21.070 3.285 21.410 3.620 ;
        RECT 25.550 3.285 25.890 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 28.990 4.350 ;
        RECT -0.430 1.760 9.450 1.885 ;
        RECT 27.395 1.760 28.990 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 28.990 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 0.635 ;
        RECT 2.430 0.300 2.770 0.635 ;
        RECT 4.670 0.300 5.010 0.635 ;
        RECT 6.910 0.300 7.250 0.635 ;
        RECT 9.150 0.300 9.490 0.635 ;
        RECT 0.000 -0.300 28.560 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 9.265 1.095 18.050 1.220 ;
        RECT 1.310 0.990 18.050 1.095 ;
        RECT 1.310 0.865 9.495 0.990 ;
        RECT 9.860 0.530 28.360 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai222_4
MACRO gf180mcu_fd_sc_mcu7t5v0__or2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.660 1.075 1.080 2.880 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.780 1.740 2.140 3.345 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 3.500 2.290 4.130 3.345 ;
        RECT 3.800 1.040 4.130 2.290 ;
        RECT 3.365 0.610 4.130 1.040 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 4.480 4.220 ;
        RECT 2.780 2.530 3.010 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 4.910 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 0.300 0.530 0.825 ;
        RECT 2.780 0.300 3.010 0.850 ;
        RECT 0.000 -0.300 4.480 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.335 3.130 1.540 3.360 ;
        RECT 1.310 1.510 1.540 3.130 ;
        RECT 2.680 1.510 3.535 1.640 ;
        RECT 1.310 1.280 3.535 1.510 ;
        RECT 1.310 0.530 1.705 1.280 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or2_1
MACRO gf180mcu_fd_sc_mcu7t5v0__or2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.660 1.015 1.020 2.280 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.780 1.430 2.140 3.390 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.121800 ;
    PORT
      LAYER Metal1 ;
        RECT 3.480 0.530 3.835 3.390 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.600 4.220 ;
        RECT 2.435 2.530 2.665 3.620 ;
        RECT 4.625 2.530 4.855 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 6.030 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 0.635 ;
        RECT 2.430 0.300 2.770 0.635 ;
        RECT 4.725 0.300 4.955 1.045 ;
        RECT 0.000 -0.300 5.600 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 2.765 0.575 3.390 ;
        RECT 0.345 2.530 1.530 2.765 ;
        RECT 1.300 1.115 1.530 2.530 ;
        RECT 2.975 1.115 3.205 2.115 ;
        RECT 1.300 0.885 3.205 1.115 ;
        RECT 1.300 0.530 1.595 0.885 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or2_2
MACRO gf180mcu_fd_sc_mcu7t5v0__or2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.595 1.800 3.500 2.120 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.870 2.360 4.275 2.680 ;
        RECT 0.870 1.765 1.210 2.360 ;
        RECT 3.930 1.825 4.275 2.360 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.304600 ;
    PORT
      LAYER Metal1 ;
        RECT 6.085 2.680 6.315 3.390 ;
        RECT 8.175 2.680 8.405 3.390 ;
        RECT 6.085 2.360 9.460 2.680 ;
        RECT 9.205 1.540 9.460 2.360 ;
        RECT 5.985 1.265 9.460 1.540 ;
        RECT 5.985 1.260 8.455 1.265 ;
        RECT 5.985 0.530 6.215 1.260 ;
        RECT 8.225 0.530 8.455 1.260 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 10.080 4.220 ;
        RECT 0.345 2.530 0.575 3.620 ;
        RECT 4.965 2.530 5.195 3.620 ;
        RECT 7.105 2.935 7.335 3.620 ;
        RECT 9.245 2.940 9.475 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 10.510 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.070 ;
        RECT 2.485 0.300 2.715 1.070 ;
        RECT 4.725 0.300 4.955 1.070 ;
        RECT 7.105 0.300 7.335 0.985 ;
        RECT 9.345 0.300 9.575 0.980 ;
        RECT 0.000 -0.300 10.080 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 2.350 2.945 4.735 3.215 ;
        RECT 4.505 2.095 4.735 2.945 ;
        RECT 4.505 1.825 8.960 2.095 ;
        RECT 4.505 1.570 4.735 1.825 ;
        RECT 1.365 1.325 4.735 1.570 ;
        RECT 1.365 0.530 1.595 1.325 ;
        RECT 3.605 0.530 3.835 1.325 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or2_4
MACRO gf180mcu_fd_sc_mcu7t5v0__or3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.520000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.660 1.595 1.020 2.855 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.520000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.780 1.595 2.140 3.390 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.520000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.900 1.595 3.350 3.390 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 4.985 0.530 5.455 3.390 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.600 4.220 ;
        RECT 3.965 2.530 4.195 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 6.030 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.310 0.300 1.650 0.735 ;
        RECT 3.730 0.300 4.070 0.735 ;
        RECT 0.000 -0.300 5.600 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.180 3.160 1.515 3.390 ;
        RECT 1.285 1.200 1.515 3.160 ;
        RECT 4.445 1.200 4.675 2.220 ;
        RECT 0.190 0.965 4.675 1.200 ;
        RECT 0.190 0.530 0.530 0.965 ;
        RECT 2.430 0.530 2.770 0.965 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or3_1
MACRO gf180mcu_fd_sc_mcu7t5v0__or3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.009000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.220 2.140 1.560 3.380 ;
        RECT 0.840 1.730 1.560 2.140 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.009000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.790 1.610 2.140 3.380 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.009000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.900 1.610 3.260 3.380 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal1 ;
        RECT 4.840 2.655 5.460 3.380 ;
        RECT 4.840 2.380 6.040 2.655 ;
        RECT 5.745 1.535 6.040 2.380 ;
        RECT 4.870 1.265 6.040 1.535 ;
        RECT 4.870 0.530 5.490 1.265 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 6.720 4.220 ;
        RECT 3.715 2.530 3.945 3.620 ;
        RECT 5.925 2.935 6.155 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 7.150 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.150 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 0.895 ;
        RECT 3.605 0.300 3.835 0.895 ;
        RECT 6.025 0.300 6.255 0.920 ;
        RECT 0.000 -0.300 6.720 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.245 1.360 0.575 3.390 ;
        RECT 3.960 1.765 5.515 1.995 ;
        RECT 3.960 1.360 4.190 1.765 ;
        RECT 0.245 1.125 4.190 1.360 ;
        RECT 0.245 0.530 0.475 1.125 ;
        RECT 2.485 0.530 2.715 1.125 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or3_2
MACRO gf180mcu_fd_sc_mcu7t5v0__or3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.320 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.910 1.325 6.105 1.590 ;
        RECT 3.495 1.170 3.785 1.325 ;
        RECT 5.735 1.170 6.105 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.530 1.820 5.550 2.105 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.870 2.380 6.175 2.655 ;
        RECT 0.870 1.820 1.160 2.380 ;
        RECT 5.945 2.115 6.175 2.380 ;
        RECT 5.945 1.820 6.570 2.115 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.243600 ;
    PORT
      LAYER Metal1 ;
        RECT 8.315 2.680 8.545 3.390 ;
        RECT 10.455 2.680 10.685 3.390 ;
        RECT 8.315 2.360 11.620 2.680 ;
        RECT 11.345 1.535 11.620 2.360 ;
        RECT 8.265 1.265 11.620 1.535 ;
        RECT 8.265 0.530 8.495 1.265 ;
        RECT 10.505 0.530 10.735 1.265 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 12.320 4.220 ;
        RECT 0.345 2.530 0.575 3.620 ;
        RECT 6.865 3.060 7.095 3.620 ;
        RECT 9.335 3.000 9.565 3.620 ;
        RECT 11.525 3.000 11.755 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 12.750 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.750 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.005 ;
        RECT 2.430 0.300 2.770 0.635 ;
        RECT 4.670 0.300 5.010 0.635 ;
        RECT 6.910 0.300 7.250 0.635 ;
        RECT 9.385 0.300 9.615 0.900 ;
        RECT 11.625 0.300 11.855 0.970 ;
        RECT 0.000 -0.300 12.320 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.505 2.935 6.635 3.220 ;
        RECT 6.405 2.755 6.635 2.935 ;
        RECT 6.405 2.520 7.030 2.755 ;
        RECT 6.800 1.995 7.030 2.520 ;
        RECT 6.800 1.765 11.095 1.995 ;
        RECT 6.800 1.095 7.030 1.765 ;
        RECT 1.940 0.920 3.260 1.095 ;
        RECT 4.190 0.920 5.495 1.095 ;
        RECT 6.360 0.920 7.030 1.095 ;
        RECT 1.940 0.865 7.030 0.920 ;
        RECT 1.940 0.775 2.185 0.865 ;
        RECT 1.265 0.545 2.185 0.775 ;
        RECT 3.015 0.545 4.430 0.865 ;
        RECT 5.260 0.545 6.620 0.865 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or3_4
MACRO gf180mcu_fd_sc_mcu7t5v0__or4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.660 1.085 1.020 2.870 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.780 1.580 2.260 3.280 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.900 1.580 3.380 3.280 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.496000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.020 1.580 4.500 3.280 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 6.070 0.630 6.575 3.380 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 6.720 4.220 ;
        RECT 5.085 2.530 5.315 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 7.150 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.150 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 0.760 ;
        RECT 2.610 0.300 2.950 0.760 ;
        RECT 5.085 0.300 5.315 0.855 ;
        RECT 0.000 -0.300 6.720 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.280 3.120 1.530 3.350 ;
        RECT 1.300 1.330 1.530 3.120 ;
        RECT 5.515 1.330 5.765 2.270 ;
        RECT 1.300 1.095 5.765 1.330 ;
        RECT 1.490 0.530 1.830 1.095 ;
        RECT 3.730 0.530 4.070 1.095 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or4_1
MACRO gf180mcu_fd_sc_mcu7t5v0__or4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.889000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.660 1.015 1.020 2.290 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.889000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.780 1.480 2.140 3.390 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.889000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.900 1.480 3.260 3.390 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.889000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.020 1.480 4.380 3.390 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.121800 ;
    PORT
      LAYER Metal1 ;
        RECT 5.970 2.680 6.585 3.390 ;
        RECT 5.970 2.360 7.280 2.680 ;
        RECT 7.010 1.560 7.280 2.360 ;
        RECT 6.025 1.240 7.280 1.560 ;
        RECT 6.025 0.530 6.585 1.240 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.840 4.220 ;
        RECT 4.820 2.530 5.050 3.620 ;
        RECT 7.045 2.990 7.275 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 8.270 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 0.655 ;
        RECT 2.430 0.300 2.770 0.655 ;
        RECT 4.670 0.300 5.010 0.655 ;
        RECT 7.145 0.300 7.375 0.900 ;
        RECT 0.000 -0.300 7.840 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 2.760 0.575 3.390 ;
        RECT 0.345 2.530 1.540 2.760 ;
        RECT 1.310 1.180 1.540 2.530 ;
        RECT 5.030 1.845 6.750 2.075 ;
        RECT 5.030 1.180 5.260 1.845 ;
        RECT 1.310 0.945 5.260 1.180 ;
        RECT 1.310 0.530 1.650 0.945 ;
        RECT 3.550 0.530 3.890 0.945 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or4_2
MACRO gf180mcu_fd_sc_mcu7t5v0__or4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.405 1.205 4.025 1.545 ;
        RECT 5.645 1.205 6.275 1.545 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.330 2.010 3.535 2.120 ;
        RECT 2.330 1.780 6.730 2.010 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.785 2.470 3.980 2.680 ;
        RECT 1.785 2.360 7.720 2.470 ;
        RECT 1.785 1.575 2.100 2.360 ;
        RECT 3.765 2.240 7.720 2.360 ;
        RECT 7.410 1.665 7.720 2.240 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.778000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.870 2.930 4.440 3.240 ;
        RECT 0.870 2.920 8.310 2.930 ;
        RECT 0.870 1.765 1.210 2.920 ;
        RECT 4.210 2.700 8.310 2.920 ;
        RECT 7.960 1.630 8.310 2.700 ;
        RECT 7.960 1.400 8.885 1.630 ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.304600 ;
    PORT
      LAYER Metal1 ;
        RECT 10.490 2.680 10.750 3.380 ;
        RECT 12.645 2.680 12.875 3.380 ;
        RECT 10.490 2.360 13.970 2.680 ;
        RECT 13.730 1.560 13.970 2.360 ;
        RECT 10.505 1.240 13.970 1.560 ;
        RECT 10.505 0.615 10.735 1.240 ;
        RECT 12.745 0.615 12.975 1.240 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 14.560 4.220 ;
        RECT 0.345 2.555 0.575 3.620 ;
        RECT 9.380 2.530 9.610 3.620 ;
        RECT 11.575 3.040 11.805 3.620 ;
        RECT 13.765 3.040 13.995 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 14.990 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 0.655 ;
        RECT 2.485 0.300 2.715 0.710 ;
        RECT 4.725 0.300 4.955 0.710 ;
        RECT 6.965 0.300 7.195 0.710 ;
        RECT 9.150 0.300 9.490 0.655 ;
        RECT 11.625 0.300 11.855 0.830 ;
        RECT 13.865 0.300 14.095 0.830 ;
        RECT 0.000 -0.300 14.560 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 4.670 3.160 9.040 3.390 ;
        RECT 8.780 2.130 9.040 3.160 ;
        RECT 8.780 1.880 13.470 2.130 ;
        RECT 9.195 1.790 13.470 1.880 ;
        RECT 9.195 1.170 9.425 1.790 ;
        RECT 1.310 0.940 3.175 1.170 ;
        RECT 1.310 0.530 1.650 0.940 ;
        RECT 2.945 0.760 3.175 0.940 ;
        RECT 4.260 0.940 5.415 1.170 ;
        RECT 4.260 0.760 4.490 0.940 ;
        RECT 2.945 0.530 4.490 0.760 ;
        RECT 5.185 0.760 5.415 0.940 ;
        RECT 6.505 0.940 9.425 1.170 ;
        RECT 6.505 0.760 6.735 0.940 ;
        RECT 5.185 0.530 6.735 0.760 ;
        RECT 8.030 0.530 8.370 0.940 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or4_4
MACRO gf180mcu_fd_sc_mcu7t5v0__sdffq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.280 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.410 1.795 5.085 2.215 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 0.595 1.030 2.150 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.825 0.595 2.150 2.150 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.739000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.465 1.795 6.630 2.200 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.893200 ;
    PORT
      LAYER Metal1 ;
        RECT 20.790 0.615 21.150 3.365 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 21.280 4.220 ;
        RECT 1.260 2.845 1.600 3.620 ;
        RECT 5.250 3.180 5.590 3.620 ;
        RECT 7.570 3.350 7.910 3.620 ;
        RECT 12.930 2.995 13.270 3.620 ;
        RECT 17.250 2.845 17.590 3.620 ;
        RECT 19.735 2.460 19.965 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 21.710 4.350 ;
        RECT -0.430 1.760 6.245 1.885 ;
        RECT 10.000 1.760 21.710 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 6.245 1.760 10.000 1.885 ;
        RECT -0.430 -0.430 21.710 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 1.140 ;
        RECT 5.295 0.300 5.635 1.075 ;
        RECT 7.780 0.300 8.010 1.045 ;
        RECT 12.980 0.300 13.320 1.085 ;
        RECT 17.625 0.300 17.855 0.680 ;
        RECT 19.685 0.300 19.915 0.995 ;
        RECT 0.000 -0.300 21.280 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 5.875 3.120 7.320 3.320 ;
        RECT 8.370 3.120 10.015 3.350 ;
        RECT 5.875 3.090 8.600 3.120 ;
        RECT 0.245 2.615 0.475 3.015 ;
        RECT 5.875 2.935 6.105 3.090 ;
        RECT 3.030 2.705 6.105 2.935 ;
        RECT 7.090 2.890 8.600 3.090 ;
        RECT 6.585 2.660 6.815 2.860 ;
        RECT 0.245 2.385 2.775 2.615 ;
        RECT 6.585 2.430 8.600 2.660 ;
        RECT 0.245 0.790 0.475 2.385 ;
        RECT 2.545 1.625 2.775 2.385 ;
        RECT 4.425 1.305 6.320 1.535 ;
        RECT 4.425 1.075 4.655 1.305 ;
        RECT 3.270 0.845 4.655 1.075 ;
        RECT 6.090 0.760 6.320 1.305 ;
        RECT 6.860 1.275 7.090 2.430 ;
        RECT 8.370 1.875 8.600 2.430 ;
        RECT 8.900 2.050 9.130 2.860 ;
        RECT 9.785 2.690 10.015 3.120 ;
        RECT 10.325 3.150 12.490 3.390 ;
        RECT 10.325 2.050 10.555 3.150 ;
        RECT 8.900 1.820 10.555 2.050 ;
        RECT 6.750 0.990 7.090 1.275 ;
        RECT 7.320 1.305 8.605 1.535 ;
        RECT 7.320 0.760 7.550 1.305 ;
        RECT 6.090 0.530 7.550 0.760 ;
        RECT 8.375 0.760 8.605 1.305 ;
        RECT 9.065 1.275 9.295 1.820 ;
        RECT 10.855 1.700 11.085 2.870 ;
        RECT 12.260 2.765 12.490 3.150 ;
        RECT 13.670 3.160 16.245 3.390 ;
        RECT 13.670 2.765 13.900 3.160 ;
        RECT 12.260 2.530 13.900 2.765 ;
        RECT 14.325 2.300 14.555 2.870 ;
        RECT 12.200 2.070 14.555 2.300 ;
        RECT 10.855 1.470 13.965 1.700 ;
        RECT 9.065 0.990 9.405 1.275 ;
        RECT 9.840 0.760 10.070 1.140 ;
        RECT 10.960 0.800 11.190 1.470 ;
        RECT 14.325 0.800 14.555 2.070 ;
        RECT 14.785 1.260 15.015 3.160 ;
        RECT 15.445 1.775 15.675 2.870 ;
        RECT 15.905 2.070 16.245 3.160 ;
        RECT 16.505 2.315 18.170 2.550 ;
        RECT 16.505 1.775 16.735 2.315 ;
        RECT 15.445 1.540 16.735 1.775 ;
        RECT 17.830 1.670 18.170 2.315 ;
        RECT 18.465 2.010 18.695 2.950 ;
        RECT 18.465 1.780 20.540 2.010 ;
        RECT 15.445 0.800 15.675 1.540 ;
        RECT 16.965 1.230 17.195 1.600 ;
        RECT 18.965 1.230 19.195 1.780 ;
        RECT 16.965 0.995 19.195 1.230 ;
        RECT 18.965 0.760 19.195 0.995 ;
        RECT 8.375 0.530 10.070 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffq_1
MACRO gf180mcu_fd_sc_mcu7t5v0__sdffq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.400 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.410 1.795 5.140 2.215 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 0.595 1.030 2.150 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.825 0.595 2.150 2.150 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.739000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.465 1.795 6.630 2.200 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.116350 ;
    PORT
      LAYER Metal1 ;
        RECT 20.760 0.615 21.180 3.390 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 22.400 4.220 ;
        RECT 1.260 2.845 1.600 3.620 ;
        RECT 5.250 3.180 5.590 3.620 ;
        RECT 7.570 3.350 7.910 3.620 ;
        RECT 12.930 2.995 13.270 3.620 ;
        RECT 17.710 2.800 18.050 3.620 ;
        RECT 19.785 2.460 20.015 3.620 ;
        RECT 21.875 2.460 22.105 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 22.830 4.350 ;
        RECT -0.430 1.760 6.245 1.885 ;
        RECT 10.000 1.760 22.830 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 6.245 1.760 10.000 1.885 ;
        RECT -0.430 -0.430 22.830 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 1.140 ;
        RECT 5.295 0.300 5.635 1.075 ;
        RECT 7.780 0.300 8.010 1.045 ;
        RECT 12.980 0.300 13.320 1.085 ;
        RECT 17.845 0.300 18.075 0.725 ;
        RECT 19.685 0.300 19.915 0.950 ;
        RECT 21.925 0.300 22.155 0.950 ;
        RECT 0.000 -0.300 22.400 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 5.875 3.120 7.320 3.320 ;
        RECT 8.370 3.120 10.015 3.350 ;
        RECT 5.875 3.090 8.600 3.120 ;
        RECT 0.245 2.615 0.475 3.015 ;
        RECT 5.875 2.935 6.105 3.090 ;
        RECT 3.030 2.705 6.105 2.935 ;
        RECT 7.090 2.890 8.600 3.090 ;
        RECT 6.585 2.660 6.815 2.860 ;
        RECT 0.245 2.385 2.775 2.615 ;
        RECT 6.585 2.430 8.600 2.660 ;
        RECT 0.245 0.790 0.475 2.385 ;
        RECT 2.545 1.625 2.775 2.385 ;
        RECT 4.425 1.305 6.265 1.535 ;
        RECT 4.425 1.075 4.655 1.305 ;
        RECT 3.270 0.845 4.655 1.075 ;
        RECT 6.035 0.760 6.265 1.305 ;
        RECT 6.860 1.275 7.090 2.430 ;
        RECT 8.370 1.875 8.600 2.430 ;
        RECT 8.900 2.050 9.130 2.860 ;
        RECT 9.785 2.690 10.015 3.120 ;
        RECT 10.325 3.150 12.490 3.390 ;
        RECT 10.325 2.050 10.555 3.150 ;
        RECT 8.900 1.820 10.555 2.050 ;
        RECT 6.750 0.990 7.090 1.275 ;
        RECT 7.320 1.305 8.605 1.535 ;
        RECT 7.320 0.760 7.550 1.305 ;
        RECT 6.035 0.530 7.550 0.760 ;
        RECT 8.375 0.760 8.605 1.305 ;
        RECT 9.065 1.275 9.295 1.820 ;
        RECT 10.855 1.700 11.085 2.870 ;
        RECT 12.260 2.765 12.490 3.150 ;
        RECT 13.670 3.160 16.245 3.390 ;
        RECT 13.670 2.765 13.900 3.160 ;
        RECT 12.260 2.530 13.900 2.765 ;
        RECT 14.325 2.300 14.555 2.870 ;
        RECT 12.200 2.070 14.555 2.300 ;
        RECT 10.855 1.470 13.965 1.700 ;
        RECT 9.065 0.990 9.405 1.275 ;
        RECT 9.840 0.760 10.070 1.140 ;
        RECT 10.960 0.800 11.190 1.470 ;
        RECT 14.285 0.800 14.555 2.070 ;
        RECT 14.785 1.260 15.015 3.160 ;
        RECT 15.425 1.775 15.675 2.870 ;
        RECT 15.905 2.070 16.245 3.160 ;
        RECT 16.655 2.315 18.630 2.550 ;
        RECT 16.655 1.775 16.885 2.315 ;
        RECT 15.425 1.540 16.885 1.775 ;
        RECT 15.425 0.800 15.675 1.540 ;
        RECT 17.200 1.230 17.450 2.080 ;
        RECT 18.290 1.460 18.630 2.315 ;
        RECT 18.965 1.795 19.195 3.345 ;
        RECT 20.245 1.795 20.515 2.085 ;
        RECT 18.965 1.565 20.515 1.795 ;
        RECT 18.965 1.230 19.195 1.565 ;
        RECT 20.245 1.275 20.515 1.565 ;
        RECT 17.200 0.995 19.195 1.230 ;
        RECT 8.375 0.530 10.070 0.760 ;
        RECT 18.965 0.575 19.195 0.995 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffq_2
MACRO gf180mcu_fd_sc_mcu7t5v0__sdffq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.640 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.410 1.795 5.180 2.215 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 0.600 1.030 2.155 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.825 0.600 2.150 2.155 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.739000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.465 1.795 6.630 2.190 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.232700 ;
    PORT
      LAYER Metal1 ;
        RECT 20.760 2.160 21.180 3.390 ;
        RECT 22.980 2.160 23.400 3.390 ;
        RECT 20.760 1.740 23.400 2.160 ;
        RECT 20.760 0.615 21.180 1.740 ;
        RECT 22.980 0.615 23.400 1.740 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 24.640 4.220 ;
        RECT 1.260 2.845 1.600 3.620 ;
        RECT 5.250 3.180 5.590 3.620 ;
        RECT 7.570 3.350 7.910 3.620 ;
        RECT 12.930 2.995 13.270 3.620 ;
        RECT 17.710 2.800 18.050 3.620 ;
        RECT 19.785 2.460 20.015 3.620 ;
        RECT 21.945 2.460 22.175 3.620 ;
        RECT 24.115 2.460 24.345 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 25.070 4.350 ;
        RECT -0.430 1.760 6.245 1.885 ;
        RECT 10.000 1.760 25.070 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 6.245 1.760 10.000 1.885 ;
        RECT -0.430 -0.430 25.070 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 1.140 ;
        RECT 5.295 0.300 5.635 1.075 ;
        RECT 7.780 0.300 8.010 1.045 ;
        RECT 12.980 0.300 13.320 1.085 ;
        RECT 17.845 0.300 18.075 0.725 ;
        RECT 19.685 0.300 19.915 0.950 ;
        RECT 21.925 0.300 22.155 0.950 ;
        RECT 24.165 0.300 24.395 0.950 ;
        RECT 0.000 -0.300 24.640 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 5.875 3.120 7.320 3.320 ;
        RECT 8.370 3.120 10.015 3.350 ;
        RECT 5.875 3.090 8.600 3.120 ;
        RECT 0.245 2.615 0.475 3.015 ;
        RECT 5.875 2.935 6.105 3.090 ;
        RECT 3.030 2.705 6.105 2.935 ;
        RECT 7.090 2.890 8.600 3.090 ;
        RECT 6.585 2.660 6.815 2.860 ;
        RECT 0.245 2.385 2.775 2.615 ;
        RECT 6.585 2.430 8.600 2.660 ;
        RECT 0.245 0.790 0.475 2.385 ;
        RECT 2.545 1.625 2.775 2.385 ;
        RECT 4.425 1.305 6.260 1.535 ;
        RECT 4.425 1.075 4.655 1.305 ;
        RECT 3.270 0.845 4.655 1.075 ;
        RECT 6.030 0.760 6.260 1.305 ;
        RECT 6.860 1.275 7.090 2.430 ;
        RECT 8.370 1.875 8.600 2.430 ;
        RECT 8.900 2.050 9.130 2.860 ;
        RECT 9.785 2.690 10.015 3.120 ;
        RECT 10.325 3.150 12.490 3.390 ;
        RECT 10.325 2.050 10.555 3.150 ;
        RECT 8.900 1.820 10.555 2.050 ;
        RECT 6.750 0.990 7.090 1.275 ;
        RECT 7.320 1.305 8.605 1.535 ;
        RECT 7.320 0.760 7.550 1.305 ;
        RECT 6.030 0.530 7.550 0.760 ;
        RECT 8.375 0.760 8.605 1.305 ;
        RECT 9.065 1.275 9.295 1.820 ;
        RECT 10.855 1.700 11.085 2.870 ;
        RECT 12.260 2.765 12.490 3.150 ;
        RECT 13.670 3.160 16.245 3.390 ;
        RECT 13.670 2.765 13.900 3.160 ;
        RECT 12.260 2.530 13.900 2.765 ;
        RECT 14.325 2.300 14.555 2.870 ;
        RECT 12.200 2.070 14.555 2.300 ;
        RECT 10.855 1.470 13.965 1.700 ;
        RECT 9.065 0.990 9.405 1.275 ;
        RECT 9.840 0.760 10.070 1.140 ;
        RECT 10.960 0.800 11.190 1.470 ;
        RECT 14.285 0.800 14.515 2.070 ;
        RECT 14.785 1.260 15.015 3.160 ;
        RECT 15.425 1.775 15.675 2.870 ;
        RECT 15.905 2.070 16.245 3.160 ;
        RECT 16.655 2.315 18.630 2.550 ;
        RECT 16.655 1.775 16.885 2.315 ;
        RECT 15.425 1.540 16.885 1.775 ;
        RECT 15.425 0.800 15.675 1.540 ;
        RECT 17.195 1.230 17.455 2.080 ;
        RECT 18.290 1.460 18.630 2.315 ;
        RECT 18.965 1.795 19.195 3.345 ;
        RECT 20.245 1.795 20.515 2.085 ;
        RECT 18.965 1.565 20.515 1.795 ;
        RECT 18.965 1.230 19.195 1.565 ;
        RECT 20.245 1.275 20.515 1.565 ;
        RECT 17.195 0.995 19.195 1.230 ;
        RECT 8.375 0.530 10.070 0.760 ;
        RECT 18.965 0.575 19.195 0.995 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffq_4
MACRO gf180mcu_fd_sc_mcu7t5v0__sdffrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffrnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.080 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.095 1.765 4.390 2.190 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.155 1.210 20.410 1.635 ;
        RECT 20.040 1.020 20.410 1.210 ;
        RECT 20.040 0.645 20.670 1.020 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 0.595 1.030 2.150 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.825 0.595 2.150 2.150 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.741500 ;
    PORT
      LAYER Metal1 ;
        RECT 5.130 1.765 6.630 2.155 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER Metal1 ;
        RECT 23.590 0.555 23.950 3.380 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 24.080 4.220 ;
        RECT 1.260 2.845 1.600 3.620 ;
        RECT 5.375 2.885 5.605 3.620 ;
        RECT 7.590 3.350 7.930 3.620 ;
        RECT 13.120 3.000 13.460 3.620 ;
        RECT 15.135 2.665 15.365 3.620 ;
        RECT 19.480 2.845 19.820 3.620 ;
        RECT 21.675 2.675 21.905 3.620 ;
        RECT 22.535 2.360 22.765 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 24.510 4.350 ;
        RECT -0.430 1.760 5.605 1.885 ;
        RECT 20.425 1.760 24.510 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 5.605 1.760 20.425 1.885 ;
        RECT -0.430 -0.430 24.510 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 1.140 ;
        RECT 5.550 0.300 5.780 1.025 ;
        RECT 7.865 0.300 8.095 1.045 ;
        RECT 14.370 0.300 14.710 0.915 ;
        RECT 19.360 0.300 19.700 0.915 ;
        RECT 22.485 0.300 22.715 0.925 ;
        RECT 0.000 -0.300 24.080 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 6.085 3.160 7.360 3.390 ;
        RECT 0.245 2.615 0.475 3.040 ;
        RECT 3.230 2.745 5.075 2.975 ;
        RECT 4.845 2.655 5.075 2.745 ;
        RECT 6.085 2.655 6.315 3.160 ;
        RECT 7.130 3.120 7.360 3.160 ;
        RECT 8.205 3.160 10.125 3.390 ;
        RECT 8.205 3.120 8.435 3.160 ;
        RECT 7.130 2.890 8.435 3.120 ;
        RECT 0.245 2.385 2.855 2.615 ;
        RECT 4.845 2.420 6.315 2.655 ;
        RECT 6.610 2.620 6.840 2.890 ;
        RECT 6.610 2.385 8.535 2.620 ;
        RECT 0.245 0.780 0.475 2.385 ;
        RECT 2.625 1.535 2.855 2.385 ;
        RECT 4.630 1.535 4.860 1.750 ;
        RECT 2.625 1.305 4.860 1.535 ;
        RECT 5.090 1.260 6.605 1.490 ;
        RECT 6.945 1.275 7.175 2.385 ;
        RECT 8.305 1.910 8.535 2.385 ;
        RECT 8.885 2.035 9.115 2.845 ;
        RECT 9.895 2.645 10.125 3.160 ;
        RECT 17.155 3.160 19.075 3.390 ;
        RECT 10.915 2.295 11.145 3.125 ;
        RECT 11.935 2.760 12.165 3.005 ;
        RECT 14.415 2.760 14.645 3.005 ;
        RECT 11.935 2.530 14.645 2.760 ;
        RECT 16.155 2.300 16.385 3.035 ;
        RECT 10.915 2.065 12.195 2.295 ;
        RECT 12.460 2.070 16.385 2.300 ;
        RECT 17.155 2.690 17.460 3.160 ;
        RECT 8.885 1.800 10.620 2.035 ;
        RECT 5.090 1.075 5.320 1.260 ;
        RECT 3.250 0.845 5.320 1.075 ;
        RECT 6.375 0.760 6.605 1.260 ;
        RECT 6.835 0.990 7.175 1.275 ;
        RECT 7.405 1.295 8.680 1.530 ;
        RECT 7.405 0.760 7.635 1.295 ;
        RECT 6.375 0.530 7.635 0.760 ;
        RECT 8.450 0.760 8.680 1.295 ;
        RECT 9.150 0.990 9.490 1.800 ;
        RECT 9.925 0.760 10.155 0.970 ;
        RECT 8.450 0.530 10.155 0.760 ;
        RECT 11.045 0.630 11.275 2.065 ;
        RECT 11.965 1.840 12.195 2.065 ;
        RECT 11.505 1.375 11.735 1.720 ;
        RECT 11.965 1.610 15.370 1.840 ;
        RECT 11.505 1.145 15.210 1.375 ;
        RECT 14.980 0.760 15.210 1.145 ;
        RECT 15.710 0.990 16.050 2.070 ;
        RECT 16.370 0.760 16.600 1.735 ;
        RECT 17.155 1.220 17.385 2.690 ;
        RECT 18.220 2.420 18.570 2.930 ;
        RECT 18.845 2.615 19.075 3.160 ;
        RECT 20.195 3.155 21.345 3.390 ;
        RECT 20.195 2.615 20.425 3.155 ;
        RECT 16.830 0.990 17.385 1.220 ;
        RECT 17.615 2.060 17.990 2.400 ;
        RECT 17.615 0.760 17.845 2.060 ;
        RECT 18.220 1.745 18.450 2.420 ;
        RECT 18.845 2.385 20.425 2.615 ;
        RECT 20.655 2.155 20.885 2.860 ;
        RECT 18.075 1.510 18.450 1.745 ;
        RECT 18.680 1.925 20.885 2.155 ;
        RECT 21.115 2.030 21.345 3.155 ;
        RECT 18.680 1.680 18.910 1.925 ;
        RECT 20.655 1.790 20.885 1.925 ;
        RECT 20.655 1.560 23.240 1.790 ;
        RECT 18.075 0.790 18.305 1.510 ;
        RECT 21.675 0.810 21.905 1.560 ;
        RECT 14.980 0.530 17.845 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffrnq_1
MACRO gf180mcu_fd_sc_mcu7t5v0__sdffrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffrnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.200 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.095 1.765 4.390 2.190 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.315000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.155 1.210 20.410 1.635 ;
        RECT 20.035 1.020 20.410 1.210 ;
        RECT 20.035 0.665 20.700 1.020 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 0.595 1.030 2.150 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.825 0.595 2.150 2.150 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.741500 ;
    PORT
      LAYER Metal1 ;
        RECT 5.130 1.765 6.630 2.155 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.113750 ;
    PORT
      LAYER Metal1 ;
        RECT 23.460 0.600 23.980 3.360 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 25.200 4.220 ;
        RECT 1.260 2.845 1.600 3.620 ;
        RECT 5.375 2.885 5.605 3.620 ;
        RECT 7.590 3.350 7.930 3.620 ;
        RECT 13.120 3.000 13.460 3.620 ;
        RECT 15.135 2.665 15.365 3.620 ;
        RECT 19.480 2.845 19.820 3.620 ;
        RECT 21.675 2.570 21.905 3.620 ;
        RECT 22.445 2.560 22.675 3.620 ;
        RECT 24.535 2.560 24.765 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 25.630 4.350 ;
        RECT -0.430 1.760 5.605 1.885 ;
        RECT 20.425 1.760 25.630 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 5.605 1.760 20.425 1.885 ;
        RECT -0.430 -0.430 25.630 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 1.140 ;
        RECT 5.550 0.300 5.780 1.025 ;
        RECT 7.865 0.300 8.095 1.045 ;
        RECT 14.370 0.300 14.710 0.915 ;
        RECT 19.360 0.300 19.700 0.915 ;
        RECT 22.395 0.300 22.625 0.925 ;
        RECT 24.635 0.300 24.865 0.925 ;
        RECT 0.000 -0.300 25.200 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 6.085 3.160 7.360 3.390 ;
        RECT 0.245 2.615 0.475 3.040 ;
        RECT 3.270 2.745 5.075 2.975 ;
        RECT 4.845 2.655 5.075 2.745 ;
        RECT 6.085 2.655 6.315 3.160 ;
        RECT 7.130 3.120 7.360 3.160 ;
        RECT 8.205 3.160 10.125 3.390 ;
        RECT 8.205 3.120 8.435 3.160 ;
        RECT 7.130 2.890 8.435 3.120 ;
        RECT 0.245 2.385 2.855 2.615 ;
        RECT 4.845 2.420 6.315 2.655 ;
        RECT 6.610 2.620 6.840 2.890 ;
        RECT 6.610 2.385 8.535 2.620 ;
        RECT 0.245 0.780 0.475 2.385 ;
        RECT 2.625 1.535 2.855 2.385 ;
        RECT 4.630 1.535 4.860 1.750 ;
        RECT 2.625 1.305 4.860 1.535 ;
        RECT 5.090 1.260 6.605 1.490 ;
        RECT 6.945 1.275 7.175 2.385 ;
        RECT 8.305 1.910 8.535 2.385 ;
        RECT 8.885 2.035 9.115 2.845 ;
        RECT 9.895 2.645 10.125 3.160 ;
        RECT 17.155 3.160 19.075 3.390 ;
        RECT 10.915 2.295 11.145 3.125 ;
        RECT 11.935 2.760 12.165 3.005 ;
        RECT 14.415 2.760 14.645 3.005 ;
        RECT 11.935 2.530 14.645 2.760 ;
        RECT 16.155 2.300 16.385 3.035 ;
        RECT 10.915 2.065 12.195 2.295 ;
        RECT 12.460 2.070 16.385 2.300 ;
        RECT 17.155 2.690 17.460 3.160 ;
        RECT 8.885 1.800 10.620 2.035 ;
        RECT 5.090 1.075 5.320 1.260 ;
        RECT 3.250 0.845 5.320 1.075 ;
        RECT 6.375 0.760 6.605 1.260 ;
        RECT 6.835 0.990 7.175 1.275 ;
        RECT 7.405 1.295 8.680 1.530 ;
        RECT 7.405 0.760 7.635 1.295 ;
        RECT 6.375 0.530 7.635 0.760 ;
        RECT 8.450 0.760 8.680 1.295 ;
        RECT 9.150 0.990 9.490 1.800 ;
        RECT 9.925 0.760 10.155 0.970 ;
        RECT 8.450 0.530 10.155 0.760 ;
        RECT 11.045 0.630 11.275 2.065 ;
        RECT 11.965 1.840 12.195 2.065 ;
        RECT 11.505 1.375 11.735 1.720 ;
        RECT 11.965 1.610 15.370 1.840 ;
        RECT 11.505 1.145 15.210 1.375 ;
        RECT 14.980 0.760 15.210 1.145 ;
        RECT 15.710 0.990 16.050 2.070 ;
        RECT 16.370 0.760 16.600 1.735 ;
        RECT 17.155 1.220 17.385 2.690 ;
        RECT 18.220 2.420 18.570 2.930 ;
        RECT 18.845 2.615 19.075 3.160 ;
        RECT 20.195 3.155 21.345 3.390 ;
        RECT 20.195 2.615 20.425 3.155 ;
        RECT 16.830 0.990 17.385 1.220 ;
        RECT 17.615 2.060 17.990 2.400 ;
        RECT 17.615 0.760 17.845 2.060 ;
        RECT 18.220 1.745 18.450 2.420 ;
        RECT 18.845 2.385 20.425 2.615 ;
        RECT 20.655 2.155 20.885 2.860 ;
        RECT 18.075 1.510 18.450 1.745 ;
        RECT 18.680 1.925 20.885 2.155 ;
        RECT 21.115 2.030 21.345 3.155 ;
        RECT 18.680 1.680 18.910 1.925 ;
        RECT 20.655 1.635 20.885 1.925 ;
        RECT 22.915 1.635 23.145 2.250 ;
        RECT 18.075 0.790 18.305 1.510 ;
        RECT 20.655 1.405 23.145 1.635 ;
        RECT 21.675 0.810 21.905 1.405 ;
        RECT 14.980 0.530 17.845 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffrnq_2
MACRO gf180mcu_fd_sc_mcu7t5v0__sdffrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffrnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.440 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.095 1.765 4.390 2.190 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.315000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.155 1.170 20.410 1.635 ;
        RECT 20.035 1.020 20.410 1.170 ;
        RECT 20.035 0.665 20.700 1.020 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 0.595 1.030 2.150 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.825 0.595 2.150 2.150 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.741500 ;
    PORT
      LAYER Metal1 ;
        RECT 5.090 1.765 6.630 2.155 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.227500 ;
    PORT
      LAYER Metal1 ;
        RECT 23.460 2.180 23.980 3.360 ;
        RECT 25.700 2.180 26.220 3.360 ;
        RECT 23.460 1.660 26.220 2.180 ;
        RECT 23.460 0.600 23.980 1.660 ;
        RECT 25.700 0.600 26.220 1.660 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 27.440 4.220 ;
        RECT 1.260 2.845 1.600 3.620 ;
        RECT 5.375 2.885 5.605 3.620 ;
        RECT 7.590 3.350 7.930 3.620 ;
        RECT 13.120 3.000 13.460 3.620 ;
        RECT 15.135 2.665 15.365 3.620 ;
        RECT 19.480 2.845 19.820 3.620 ;
        RECT 21.675 2.535 21.905 3.620 ;
        RECT 22.445 2.560 22.675 3.620 ;
        RECT 24.610 2.560 24.840 3.620 ;
        RECT 26.775 2.560 27.005 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 27.870 4.350 ;
        RECT -0.430 1.760 5.605 1.885 ;
        RECT 20.425 1.760 27.870 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 5.605 1.760 20.425 1.885 ;
        RECT -0.430 -0.430 27.870 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 1.140 ;
        RECT 5.550 0.300 5.780 1.025 ;
        RECT 7.865 0.300 8.095 1.045 ;
        RECT 14.370 0.300 14.710 0.915 ;
        RECT 19.360 0.300 19.700 0.915 ;
        RECT 22.395 0.300 22.625 0.925 ;
        RECT 24.635 0.300 24.865 0.925 ;
        RECT 26.875 0.300 27.105 0.925 ;
        RECT 0.000 -0.300 27.440 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 6.085 3.160 7.360 3.390 ;
        RECT 0.245 2.615 0.475 3.040 ;
        RECT 3.270 2.745 5.075 2.975 ;
        RECT 4.845 2.655 5.075 2.745 ;
        RECT 6.085 2.655 6.315 3.160 ;
        RECT 7.130 3.120 7.360 3.160 ;
        RECT 8.205 3.160 10.125 3.390 ;
        RECT 8.205 3.120 8.435 3.160 ;
        RECT 7.130 2.890 8.435 3.120 ;
        RECT 0.245 2.385 2.855 2.615 ;
        RECT 4.845 2.420 6.315 2.655 ;
        RECT 6.610 2.620 6.840 2.890 ;
        RECT 6.610 2.385 8.535 2.620 ;
        RECT 0.245 0.780 0.475 2.385 ;
        RECT 2.625 1.535 2.855 2.385 ;
        RECT 4.630 1.535 4.860 1.750 ;
        RECT 2.625 1.305 4.860 1.535 ;
        RECT 5.090 1.260 6.605 1.490 ;
        RECT 6.945 1.275 7.175 2.385 ;
        RECT 8.305 1.910 8.535 2.385 ;
        RECT 8.885 2.035 9.115 2.845 ;
        RECT 9.895 2.645 10.125 3.160 ;
        RECT 17.155 3.160 19.075 3.390 ;
        RECT 10.915 2.295 11.145 3.125 ;
        RECT 11.935 2.760 12.165 3.005 ;
        RECT 14.415 2.760 14.645 3.005 ;
        RECT 11.935 2.530 14.645 2.760 ;
        RECT 16.155 2.300 16.385 3.035 ;
        RECT 10.915 2.065 12.195 2.295 ;
        RECT 12.460 2.070 16.385 2.300 ;
        RECT 17.155 2.690 17.460 3.160 ;
        RECT 8.885 1.800 10.620 2.035 ;
        RECT 5.090 1.075 5.320 1.260 ;
        RECT 3.250 0.845 5.320 1.075 ;
        RECT 6.375 0.760 6.605 1.260 ;
        RECT 6.835 0.990 7.175 1.275 ;
        RECT 7.405 1.295 8.680 1.530 ;
        RECT 7.405 0.760 7.635 1.295 ;
        RECT 6.375 0.530 7.635 0.760 ;
        RECT 8.450 0.760 8.680 1.295 ;
        RECT 9.150 0.990 9.490 1.800 ;
        RECT 9.925 0.760 10.155 0.970 ;
        RECT 8.450 0.530 10.155 0.760 ;
        RECT 11.045 0.630 11.275 2.065 ;
        RECT 11.965 1.840 12.195 2.065 ;
        RECT 11.505 1.375 11.735 1.720 ;
        RECT 11.965 1.610 15.370 1.840 ;
        RECT 11.505 1.145 15.210 1.375 ;
        RECT 14.980 0.760 15.210 1.145 ;
        RECT 15.710 0.990 16.050 2.070 ;
        RECT 16.370 0.760 16.600 1.735 ;
        RECT 17.155 1.220 17.385 2.690 ;
        RECT 18.220 2.420 18.570 2.930 ;
        RECT 18.845 2.615 19.075 3.160 ;
        RECT 20.195 3.155 21.345 3.390 ;
        RECT 20.195 2.615 20.425 3.155 ;
        RECT 16.830 0.990 17.385 1.220 ;
        RECT 17.615 2.060 17.990 2.400 ;
        RECT 17.615 0.760 17.845 2.060 ;
        RECT 18.220 1.745 18.450 2.420 ;
        RECT 18.845 2.385 20.425 2.615 ;
        RECT 20.655 2.155 20.885 2.860 ;
        RECT 18.075 1.510 18.450 1.745 ;
        RECT 18.680 1.925 20.885 2.155 ;
        RECT 21.115 2.030 21.345 3.155 ;
        RECT 18.680 1.680 18.910 1.925 ;
        RECT 20.655 1.635 20.885 1.925 ;
        RECT 22.915 1.635 23.145 2.250 ;
        RECT 18.075 0.790 18.305 1.510 ;
        RECT 20.655 1.405 23.145 1.635 ;
        RECT 21.675 0.810 21.905 1.405 ;
        RECT 14.980 0.530 17.845 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffrnq_4
MACRO gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.880 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.405 1.765 4.390 2.190 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.204500 ;
    PORT
      LAYER Metal1 ;
        RECT 22.525 1.765 23.430 2.155 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 0.595 1.030 2.150 ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062000 ;
    PORT
      LAYER Metal1 ;
        RECT 20.605 1.210 21.140 2.195 ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.825 0.595 2.150 2.150 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.741500 ;
    PORT
      LAYER Metal1 ;
        RECT 5.130 1.765 6.630 2.155 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 25.860 2.505 26.320 3.380 ;
        RECT 25.860 2.205 26.555 2.505 ;
        RECT 26.255 1.160 26.555 2.205 ;
        RECT 25.755 0.655 26.555 1.160 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 26.880 4.220 ;
        RECT 1.260 2.845 1.600 3.620 ;
        RECT 5.375 2.885 5.605 3.620 ;
        RECT 7.590 3.350 7.930 3.620 ;
        RECT 13.010 3.445 13.350 3.620 ;
        RECT 16.200 3.445 16.560 3.620 ;
        RECT 20.465 2.915 20.695 3.620 ;
        RECT 22.630 2.970 22.970 3.620 ;
        RECT 25.055 2.530 25.285 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 27.310 4.350 ;
        RECT -0.430 1.760 6.455 1.885 ;
        RECT 9.870 1.760 13.630 1.885 ;
        RECT 19.590 1.760 27.310 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 6.455 1.760 9.870 1.885 ;
        RECT 13.630 1.760 19.590 1.885 ;
        RECT -0.430 -0.430 27.310 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 1.140 ;
        RECT 5.550 0.300 5.780 1.025 ;
        RECT 7.865 0.300 8.095 1.045 ;
        RECT 13.780 0.300 14.140 0.915 ;
        RECT 21.860 0.300 22.200 1.075 ;
        RECT 25.055 0.300 25.285 1.160 ;
        RECT 0.000 -0.300 26.880 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 6.085 3.160 7.360 3.390 ;
        RECT 0.245 2.615 0.475 3.040 ;
        RECT 3.270 2.745 5.075 2.975 ;
        RECT 4.845 2.655 5.075 2.745 ;
        RECT 6.085 2.655 6.315 3.160 ;
        RECT 7.130 3.120 7.360 3.160 ;
        RECT 8.205 3.160 9.835 3.390 ;
        RECT 11.265 3.215 12.780 3.390 ;
        RECT 13.580 3.215 15.970 3.390 ;
        RECT 16.790 3.215 18.275 3.390 ;
        RECT 11.265 3.160 18.275 3.215 ;
        RECT 8.205 3.120 8.435 3.160 ;
        RECT 7.130 2.890 8.435 3.120 ;
        RECT 0.245 2.385 2.855 2.615 ;
        RECT 4.845 2.420 6.315 2.655 ;
        RECT 6.610 2.620 6.840 2.890 ;
        RECT 6.610 2.385 8.535 2.620 ;
        RECT 0.245 0.780 0.475 2.385 ;
        RECT 2.625 1.535 2.855 2.385 ;
        RECT 4.630 1.535 4.860 1.750 ;
        RECT 2.625 1.305 4.860 1.535 ;
        RECT 5.090 1.260 6.240 1.490 ;
        RECT 6.945 1.275 7.175 2.385 ;
        RECT 8.305 1.910 8.535 2.385 ;
        RECT 8.885 2.035 9.115 2.845 ;
        RECT 9.605 2.485 9.835 3.160 ;
        RECT 12.550 2.985 13.810 3.160 ;
        RECT 15.740 2.985 17.020 3.160 ;
        RECT 10.800 2.295 11.030 2.870 ;
        RECT 11.680 2.755 12.200 2.775 ;
        RECT 14.160 2.755 14.600 2.780 ;
        RECT 11.680 2.525 14.600 2.755 ;
        RECT 14.960 2.755 15.400 2.780 ;
        RECT 17.360 2.755 17.790 2.780 ;
        RECT 14.960 2.525 17.790 2.755 ;
        RECT 10.800 2.065 15.905 2.295 ;
        RECT 8.885 1.800 10.405 2.035 ;
        RECT 5.090 1.075 5.320 1.260 ;
        RECT 3.250 0.845 5.320 1.075 ;
        RECT 6.010 0.760 6.240 1.260 ;
        RECT 6.835 0.990 7.175 1.275 ;
        RECT 7.405 1.295 8.680 1.530 ;
        RECT 7.405 0.760 7.635 1.295 ;
        RECT 6.010 0.530 7.635 0.760 ;
        RECT 8.450 0.760 8.680 1.295 ;
        RECT 9.150 0.990 9.490 1.800 ;
        RECT 9.925 0.760 10.155 0.980 ;
        RECT 8.450 0.530 10.155 0.760 ;
        RECT 11.045 0.620 11.275 2.065 ;
        RECT 16.325 1.835 16.665 2.525 ;
        RECT 18.045 2.035 18.275 3.160 ;
        RECT 18.525 3.160 20.235 3.390 ;
        RECT 11.625 1.375 11.855 1.700 ;
        RECT 12.295 1.605 16.665 1.835 ;
        RECT 18.525 1.805 18.755 3.160 ;
        RECT 19.545 2.225 19.775 2.835 ;
        RECT 20.005 2.685 20.235 3.160 ;
        RECT 20.925 3.160 22.310 3.390 ;
        RECT 20.925 2.685 21.155 3.160 ;
        RECT 20.005 2.455 21.155 2.685 ;
        RECT 11.625 1.145 14.600 1.375 ;
        RECT 14.370 0.760 14.600 1.145 ;
        RECT 16.325 0.990 16.665 1.605 ;
        RECT 16.940 0.760 17.170 1.745 ;
        RECT 17.445 1.575 18.755 1.805 ;
        RECT 18.985 1.995 20.185 2.225 ;
        RECT 21.430 2.155 21.770 2.930 ;
        RECT 22.080 2.740 22.310 3.160 ;
        RECT 23.200 3.160 24.490 3.390 ;
        RECT 23.200 2.740 23.430 3.160 ;
        RECT 22.080 2.510 23.430 2.740 ;
        RECT 17.445 0.990 17.785 1.575 ;
        RECT 18.985 1.220 19.215 1.995 ;
        RECT 18.570 0.990 19.215 1.220 ;
        RECT 19.445 0.760 19.675 1.765 ;
        RECT 14.370 0.530 19.675 0.760 ;
        RECT 19.955 0.960 20.185 1.995 ;
        RECT 21.400 1.925 21.770 2.155 ;
        RECT 21.400 0.960 21.630 1.925 ;
        RECT 22.065 1.535 22.295 2.200 ;
        RECT 23.690 1.535 24.030 2.930 ;
        RECT 24.260 2.060 24.490 3.160 ;
        RECT 24.335 1.600 25.780 1.830 ;
        RECT 24.335 1.535 24.565 1.600 ;
        RECT 22.065 1.305 24.565 1.535 ;
        RECT 19.955 0.715 21.630 0.960 ;
        RECT 24.335 0.780 24.565 1.305 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_1
MACRO gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.000 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.410 1.765 4.390 2.155 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.354500 ;
    PORT
      LAYER Metal1 ;
        RECT 22.490 1.765 23.430 2.155 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 0.595 1.030 2.150 ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062000 ;
    PORT
      LAYER Metal1 ;
        RECT 20.605 1.210 21.140 2.190 ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.825 0.595 2.150 2.150 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.741500 ;
    PORT
      LAYER Metal1 ;
        RECT 5.130 1.765 6.630 2.155 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.060800 ;
    PORT
      LAYER Metal1 ;
        RECT 25.850 2.660 26.300 3.380 ;
        RECT 25.850 2.385 27.310 2.660 ;
        RECT 27.025 1.535 27.310 2.385 ;
        RECT 25.850 1.210 27.310 1.535 ;
        RECT 25.850 0.610 26.435 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 28.000 4.220 ;
        RECT 1.260 2.845 1.600 3.620 ;
        RECT 5.375 2.885 5.605 3.620 ;
        RECT 7.590 3.350 7.930 3.620 ;
        RECT 13.010 3.445 13.350 3.620 ;
        RECT 16.200 3.445 16.560 3.620 ;
        RECT 20.465 2.915 20.695 3.620 ;
        RECT 22.630 2.970 22.970 3.620 ;
        RECT 24.885 2.530 25.115 3.620 ;
        RECT 27.055 2.940 27.285 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 28.430 4.350 ;
        RECT -0.430 1.760 6.455 1.885 ;
        RECT 9.870 1.760 13.630 1.885 ;
        RECT 19.590 1.760 28.430 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 6.455 1.760 9.870 1.885 ;
        RECT 13.630 1.760 19.590 1.885 ;
        RECT -0.430 -0.430 28.430 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 1.140 ;
        RECT 5.550 0.300 5.780 1.025 ;
        RECT 7.865 0.300 8.095 1.045 ;
        RECT 13.780 0.300 14.140 0.915 ;
        RECT 21.860 0.300 22.200 1.075 ;
        RECT 25.055 0.300 25.285 0.850 ;
        RECT 27.295 0.300 27.525 0.850 ;
        RECT 0.000 -0.300 28.000 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 6.085 3.160 7.360 3.390 ;
        RECT 0.245 2.615 0.475 3.040 ;
        RECT 3.270 2.745 4.120 2.975 ;
        RECT 3.890 2.655 4.120 2.745 ;
        RECT 6.085 2.655 6.315 3.160 ;
        RECT 7.130 3.120 7.360 3.160 ;
        RECT 8.205 3.160 9.835 3.390 ;
        RECT 11.265 3.215 12.780 3.390 ;
        RECT 13.580 3.215 15.970 3.390 ;
        RECT 16.790 3.215 18.275 3.390 ;
        RECT 11.265 3.160 18.275 3.215 ;
        RECT 8.205 3.120 8.435 3.160 ;
        RECT 7.130 2.890 8.435 3.120 ;
        RECT 0.245 2.385 2.855 2.615 ;
        RECT 3.890 2.420 6.315 2.655 ;
        RECT 6.610 2.620 6.840 2.890 ;
        RECT 6.610 2.385 8.535 2.620 ;
        RECT 0.245 0.780 0.475 2.385 ;
        RECT 2.625 1.535 2.855 2.385 ;
        RECT 4.630 1.535 4.860 1.750 ;
        RECT 2.625 1.305 4.860 1.535 ;
        RECT 5.090 1.260 6.240 1.490 ;
        RECT 6.945 1.275 7.175 2.385 ;
        RECT 8.305 1.910 8.535 2.385 ;
        RECT 8.885 2.035 9.115 2.890 ;
        RECT 9.605 2.485 9.835 3.160 ;
        RECT 12.550 2.985 13.810 3.160 ;
        RECT 15.740 2.985 17.020 3.160 ;
        RECT 10.800 2.295 11.030 2.870 ;
        RECT 11.680 2.755 12.200 2.775 ;
        RECT 14.160 2.755 14.600 2.780 ;
        RECT 11.680 2.525 14.600 2.755 ;
        RECT 14.960 2.755 15.400 2.780 ;
        RECT 17.360 2.755 17.790 2.780 ;
        RECT 14.960 2.525 17.790 2.755 ;
        RECT 10.800 2.065 15.905 2.295 ;
        RECT 8.885 1.800 10.390 2.035 ;
        RECT 5.090 1.075 5.320 1.260 ;
        RECT 3.250 0.845 5.320 1.075 ;
        RECT 6.010 0.760 6.240 1.260 ;
        RECT 6.835 0.990 7.175 1.275 ;
        RECT 7.405 1.295 8.680 1.530 ;
        RECT 7.405 0.760 7.635 1.295 ;
        RECT 6.010 0.530 7.635 0.760 ;
        RECT 8.450 0.760 8.680 1.295 ;
        RECT 9.150 0.990 9.490 1.800 ;
        RECT 9.925 0.760 10.155 0.980 ;
        RECT 8.450 0.530 10.155 0.760 ;
        RECT 11.045 0.620 11.275 2.065 ;
        RECT 16.325 1.835 16.665 2.525 ;
        RECT 18.045 2.035 18.275 3.160 ;
        RECT 18.525 3.160 20.235 3.390 ;
        RECT 11.625 1.375 11.855 1.700 ;
        RECT 12.295 1.605 16.665 1.835 ;
        RECT 18.525 1.805 18.755 3.160 ;
        RECT 19.545 2.225 19.775 2.835 ;
        RECT 20.005 2.685 20.235 3.160 ;
        RECT 20.925 3.160 22.315 3.390 ;
        RECT 20.925 2.685 21.155 3.160 ;
        RECT 20.005 2.455 21.155 2.685 ;
        RECT 11.625 1.145 14.600 1.375 ;
        RECT 14.370 0.760 14.600 1.145 ;
        RECT 16.325 0.990 16.665 1.605 ;
        RECT 16.940 0.760 17.170 1.745 ;
        RECT 17.445 1.575 18.755 1.805 ;
        RECT 18.985 1.995 20.185 2.225 ;
        RECT 21.430 2.155 21.770 2.930 ;
        RECT 22.080 2.740 22.315 3.160 ;
        RECT 23.200 3.160 24.490 3.390 ;
        RECT 23.200 2.740 23.430 3.160 ;
        RECT 22.080 2.510 23.430 2.740 ;
        RECT 17.445 0.990 17.785 1.575 ;
        RECT 18.985 1.220 19.215 1.995 ;
        RECT 18.570 0.990 19.215 1.220 ;
        RECT 19.445 0.760 19.675 1.765 ;
        RECT 14.370 0.530 19.675 0.760 ;
        RECT 19.955 0.960 20.185 1.995 ;
        RECT 21.400 1.925 21.770 2.155 ;
        RECT 21.400 0.960 21.630 1.925 ;
        RECT 22.010 1.535 22.240 2.200 ;
        RECT 23.690 1.535 24.030 2.930 ;
        RECT 24.260 1.910 24.490 3.160 ;
        RECT 24.945 1.825 26.790 2.095 ;
        RECT 24.945 1.535 25.175 1.825 ;
        RECT 22.010 1.305 25.175 1.535 ;
        RECT 19.955 0.715 21.630 0.960 ;
        RECT 24.335 0.640 24.565 1.305 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_2
MACRO gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.240 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.410 1.765 4.390 2.155 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.354500 ;
    PORT
      LAYER Metal1 ;
        RECT 22.490 1.765 23.430 2.155 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 0.595 1.030 2.150 ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062000 ;
    PORT
      LAYER Metal1 ;
        RECT 20.605 1.210 21.140 2.190 ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.825 0.595 2.150 2.150 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.741500 ;
    PORT
      LAYER Metal1 ;
        RECT 5.130 1.765 6.630 2.155 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.121600 ;
    PORT
      LAYER Metal1 ;
        RECT 25.785 2.655 26.180 3.380 ;
        RECT 27.585 2.655 28.085 3.380 ;
        RECT 25.785 2.385 29.540 2.655 ;
        RECT 29.255 1.535 29.540 2.385 ;
        RECT 25.850 1.205 29.540 1.535 ;
        RECT 25.850 0.610 26.435 1.205 ;
        RECT 28.135 0.610 28.695 1.205 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 30.240 4.220 ;
        RECT 1.260 2.845 1.600 3.620 ;
        RECT 5.375 2.885 5.605 3.620 ;
        RECT 7.590 3.350 7.930 3.620 ;
        RECT 13.010 3.445 13.350 3.620 ;
        RECT 16.200 3.445 16.560 3.620 ;
        RECT 20.465 2.915 20.695 3.620 ;
        RECT 22.630 2.970 22.970 3.620 ;
        RECT 24.765 2.530 24.995 3.620 ;
        RECT 26.805 3.000 27.035 3.620 ;
        RECT 28.845 3.000 29.075 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 30.670 4.350 ;
        RECT -0.430 1.760 6.455 1.885 ;
        RECT 9.870 1.760 13.630 1.885 ;
        RECT 19.590 1.760 30.670 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 6.455 1.760 9.870 1.885 ;
        RECT 13.630 1.760 19.590 1.885 ;
        RECT -0.430 -0.430 30.670 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 1.140 ;
        RECT 5.550 0.300 5.780 1.025 ;
        RECT 7.865 0.300 8.095 1.045 ;
        RECT 13.780 0.300 14.140 0.915 ;
        RECT 21.860 0.300 22.200 1.075 ;
        RECT 25.055 0.300 25.285 0.925 ;
        RECT 27.295 0.300 27.525 0.925 ;
        RECT 29.535 0.300 29.765 0.925 ;
        RECT 0.000 -0.300 30.240 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 6.085 3.160 7.360 3.390 ;
        RECT 0.245 2.615 0.475 3.040 ;
        RECT 3.270 2.745 4.120 2.975 ;
        RECT 3.890 2.655 4.120 2.745 ;
        RECT 6.085 2.655 6.315 3.160 ;
        RECT 7.130 3.120 7.360 3.160 ;
        RECT 8.205 3.160 9.835 3.390 ;
        RECT 11.265 3.215 12.780 3.390 ;
        RECT 13.580 3.215 15.970 3.390 ;
        RECT 16.790 3.215 18.275 3.390 ;
        RECT 11.265 3.160 18.275 3.215 ;
        RECT 8.205 3.120 8.435 3.160 ;
        RECT 7.130 2.890 8.435 3.120 ;
        RECT 0.245 2.385 2.855 2.615 ;
        RECT 3.890 2.420 6.315 2.655 ;
        RECT 6.610 2.620 6.840 2.890 ;
        RECT 6.610 2.385 8.535 2.620 ;
        RECT 0.245 0.780 0.475 2.385 ;
        RECT 2.625 1.535 2.855 2.385 ;
        RECT 4.630 1.535 4.860 1.750 ;
        RECT 2.625 1.305 4.860 1.535 ;
        RECT 5.090 1.260 6.240 1.490 ;
        RECT 6.945 1.285 7.175 2.385 ;
        RECT 8.305 1.910 8.535 2.385 ;
        RECT 8.885 2.035 9.115 2.890 ;
        RECT 9.605 2.385 9.835 3.160 ;
        RECT 12.550 2.985 13.810 3.160 ;
        RECT 15.740 2.985 17.020 3.160 ;
        RECT 10.800 2.295 11.030 2.870 ;
        RECT 11.680 2.755 12.200 2.775 ;
        RECT 14.160 2.755 14.600 2.780 ;
        RECT 11.680 2.525 14.600 2.755 ;
        RECT 14.960 2.755 15.400 2.780 ;
        RECT 17.360 2.755 17.790 2.780 ;
        RECT 14.960 2.525 17.790 2.755 ;
        RECT 10.800 2.065 15.905 2.295 ;
        RECT 8.885 1.800 10.395 2.035 ;
        RECT 5.090 1.075 5.320 1.260 ;
        RECT 3.250 0.845 5.320 1.075 ;
        RECT 6.010 0.760 6.240 1.260 ;
        RECT 6.835 0.990 7.175 1.285 ;
        RECT 7.405 1.295 8.680 1.530 ;
        RECT 7.405 0.760 7.635 1.295 ;
        RECT 6.010 0.530 7.635 0.760 ;
        RECT 8.450 0.760 8.680 1.295 ;
        RECT 9.150 0.990 9.490 1.800 ;
        RECT 9.925 0.760 10.155 0.980 ;
        RECT 8.450 0.530 10.155 0.760 ;
        RECT 11.045 0.620 11.275 2.065 ;
        RECT 16.325 1.835 16.665 2.525 ;
        RECT 18.045 2.035 18.275 3.160 ;
        RECT 18.525 3.160 20.235 3.390 ;
        RECT 11.625 1.375 11.855 1.700 ;
        RECT 12.295 1.605 16.665 1.835 ;
        RECT 18.525 1.805 18.755 3.160 ;
        RECT 19.545 2.225 19.775 2.835 ;
        RECT 20.005 2.685 20.235 3.160 ;
        RECT 20.925 3.160 22.315 3.390 ;
        RECT 20.925 2.685 21.155 3.160 ;
        RECT 20.005 2.455 21.155 2.685 ;
        RECT 11.625 1.145 14.600 1.375 ;
        RECT 14.370 0.760 14.600 1.145 ;
        RECT 16.325 0.990 16.665 1.605 ;
        RECT 16.940 0.760 17.170 1.745 ;
        RECT 17.445 1.575 18.755 1.805 ;
        RECT 18.985 1.995 20.185 2.225 ;
        RECT 21.430 2.155 21.770 2.930 ;
        RECT 22.080 2.740 22.315 3.160 ;
        RECT 23.200 3.160 24.490 3.390 ;
        RECT 23.200 2.740 23.430 3.160 ;
        RECT 22.080 2.510 23.430 2.740 ;
        RECT 17.445 0.990 17.785 1.575 ;
        RECT 18.985 1.220 19.215 1.995 ;
        RECT 18.570 0.990 19.215 1.220 ;
        RECT 19.445 0.760 19.675 1.765 ;
        RECT 14.370 0.530 19.675 0.760 ;
        RECT 19.955 0.960 20.185 1.995 ;
        RECT 21.400 1.925 21.770 2.155 ;
        RECT 21.400 0.960 21.630 1.925 ;
        RECT 22.010 1.535 22.240 2.200 ;
        RECT 23.690 1.535 24.030 2.930 ;
        RECT 24.260 1.910 24.490 3.160 ;
        RECT 24.945 1.825 28.725 2.095 ;
        RECT 24.945 1.535 25.175 1.825 ;
        RECT 22.010 1.305 25.175 1.535 ;
        RECT 19.955 0.715 21.630 0.960 ;
        RECT 24.335 0.655 24.565 1.305 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_4
MACRO gf180mcu_fd_sc_mcu7t5v0__sdffsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffsnq_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.200 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.410 1.765 4.390 2.155 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 0.595 1.030 2.150 ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.057000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.620 1.170 20.110 2.190 ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.825 0.595 2.150 2.150 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.741500 ;
    PORT
      LAYER Metal1 ;
        RECT 5.130 1.765 6.630 2.155 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 24.220 0.595 24.770 3.380 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 25.200 4.220 ;
        RECT 1.260 2.845 1.600 3.620 ;
        RECT 5.375 2.885 5.605 3.620 ;
        RECT 7.590 3.350 7.930 3.620 ;
        RECT 13.190 3.445 13.530 3.620 ;
        RECT 15.460 2.910 15.820 3.620 ;
        RECT 19.470 2.965 19.810 3.620 ;
        RECT 21.590 2.965 21.930 3.620 ;
        RECT 23.515 2.530 23.745 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 25.630 4.350 ;
        RECT -0.430 1.760 6.455 1.885 ;
        RECT 9.875 1.760 12.970 1.885 ;
        RECT 18.650 1.760 25.630 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 6.455 1.760 9.875 1.885 ;
        RECT 12.970 1.760 18.650 1.885 ;
        RECT -0.430 -0.430 25.630 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 1.140 ;
        RECT 5.550 0.300 5.780 1.025 ;
        RECT 7.865 0.300 8.095 1.045 ;
        RECT 13.120 0.300 13.480 0.915 ;
        RECT 21.475 0.300 21.705 0.890 ;
        RECT 23.315 0.300 23.545 0.905 ;
        RECT 0.000 -0.300 25.200 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 6.085 3.160 7.360 3.390 ;
        RECT 0.245 2.615 0.475 3.040 ;
        RECT 3.270 2.745 4.120 2.975 ;
        RECT 3.890 2.655 4.120 2.745 ;
        RECT 6.085 2.655 6.315 3.160 ;
        RECT 7.130 3.120 7.360 3.160 ;
        RECT 8.205 3.160 9.835 3.390 ;
        RECT 11.265 3.215 12.780 3.390 ;
        RECT 13.760 3.215 15.230 3.390 ;
        RECT 11.265 3.160 15.230 3.215 ;
        RECT 8.205 3.120 8.435 3.160 ;
        RECT 7.130 2.890 8.435 3.120 ;
        RECT 0.245 2.385 2.855 2.615 ;
        RECT 3.890 2.420 6.315 2.655 ;
        RECT 6.610 2.620 6.840 2.890 ;
        RECT 6.610 2.385 8.535 2.620 ;
        RECT 0.245 0.780 0.475 2.385 ;
        RECT 2.625 1.535 2.855 2.385 ;
        RECT 4.630 1.535 4.860 1.740 ;
        RECT 2.625 1.305 4.860 1.535 ;
        RECT 5.090 1.260 6.240 1.490 ;
        RECT 6.945 1.275 7.175 2.385 ;
        RECT 8.305 1.910 8.535 2.385 ;
        RECT 8.885 2.035 9.115 2.890 ;
        RECT 9.605 2.485 9.835 3.160 ;
        RECT 12.550 2.985 13.990 3.160 ;
        RECT 10.800 2.295 11.030 2.870 ;
        RECT 10.800 2.065 14.255 2.295 ;
        RECT 14.485 2.220 14.715 2.930 ;
        RECT 15.000 2.680 15.230 3.160 ;
        RECT 16.050 3.115 17.250 3.345 ;
        RECT 16.050 2.680 16.280 3.115 ;
        RECT 15.000 2.450 16.280 2.680 ;
        RECT 16.510 2.220 16.740 2.885 ;
        RECT 8.885 1.800 10.390 2.035 ;
        RECT 5.090 1.075 5.320 1.260 ;
        RECT 3.250 0.845 5.320 1.075 ;
        RECT 6.010 0.760 6.240 1.260 ;
        RECT 6.835 0.990 7.175 1.275 ;
        RECT 7.405 1.295 8.680 1.530 ;
        RECT 7.405 0.760 7.635 1.295 ;
        RECT 6.010 0.530 7.635 0.760 ;
        RECT 8.450 0.760 8.680 1.295 ;
        RECT 9.150 0.990 9.490 1.800 ;
        RECT 9.925 0.760 10.155 0.980 ;
        RECT 8.450 0.530 10.155 0.760 ;
        RECT 11.045 0.620 11.275 2.065 ;
        RECT 14.485 1.990 16.740 2.220 ;
        RECT 17.020 2.065 17.250 3.115 ;
        RECT 17.530 3.115 19.240 3.345 ;
        RECT 14.485 1.835 14.715 1.990 ;
        RECT 11.625 1.375 11.955 1.700 ;
        RECT 12.475 1.605 14.715 1.835 ;
        RECT 11.625 1.145 14.330 1.375 ;
        RECT 14.100 0.760 14.330 1.145 ;
        RECT 15.470 0.990 15.810 1.990 ;
        RECT 17.530 1.760 17.760 3.115 ;
        RECT 18.550 2.315 18.780 2.885 ;
        RECT 19.010 2.735 19.240 3.115 ;
        RECT 20.040 3.160 21.340 3.390 ;
        RECT 20.040 2.735 20.270 3.160 ;
        RECT 19.010 2.505 20.270 2.735 ;
        RECT 16.090 0.760 16.320 1.740 ;
        RECT 16.590 1.525 17.760 1.760 ;
        RECT 17.990 2.275 18.780 2.315 ;
        RECT 17.990 2.045 19.280 2.275 ;
        RECT 16.590 0.990 16.930 1.525 ;
        RECT 17.990 1.265 18.220 2.045 ;
        RECT 17.710 0.990 18.220 1.265 ;
        RECT 18.450 0.760 18.820 1.815 ;
        RECT 14.100 0.530 18.820 0.760 ;
        RECT 19.050 0.760 19.280 2.045 ;
        RECT 20.500 0.760 20.840 2.930 ;
        RECT 21.110 2.735 21.340 3.160 ;
        RECT 21.110 2.505 22.530 2.735 ;
        RECT 21.115 1.725 21.345 2.170 ;
        RECT 22.190 1.960 22.530 2.505 ;
        RECT 22.775 1.780 23.005 3.150 ;
        RECT 22.775 1.725 23.990 1.780 ;
        RECT 21.115 1.495 23.990 1.725 ;
        RECT 19.050 0.530 20.840 0.760 ;
        RECT 22.540 1.440 23.990 1.495 ;
        RECT 22.540 0.655 22.890 1.440 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffsnq_1
MACRO gf180mcu_fd_sc_mcu7t5v0__sdffsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffsnq_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.320 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.410 1.765 4.390 2.155 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 0.595 1.030 2.150 ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.057000 ;
    PORT
      LAYER Metal1 ;
        RECT 19.620 1.170 20.110 2.190 ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.825 0.595 2.150 2.150 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.741500 ;
    PORT
      LAYER Metal1 ;
        RECT 5.130 1.765 6.630 2.155 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.079100 ;
    PORT
      LAYER Metal1 ;
        RECT 24.555 2.655 25.100 3.380 ;
        RECT 24.555 2.380 25.795 2.655 ;
        RECT 25.530 1.535 25.795 2.380 ;
        RECT 24.170 1.265 25.795 1.535 ;
        RECT 24.170 0.610 24.695 1.265 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 26.320 4.220 ;
        RECT 1.260 2.845 1.600 3.620 ;
        RECT 5.375 2.885 5.605 3.620 ;
        RECT 7.590 3.350 7.930 3.620 ;
        RECT 13.190 3.445 13.530 3.620 ;
        RECT 15.460 2.910 15.820 3.620 ;
        RECT 19.485 2.965 19.825 3.620 ;
        RECT 21.580 2.965 21.920 3.620 ;
        RECT 23.540 2.530 23.770 3.620 ;
        RECT 25.595 2.945 25.825 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 26.750 4.350 ;
        RECT -0.430 1.760 6.455 1.885 ;
        RECT 9.870 1.760 12.970 1.885 ;
        RECT 18.650 1.760 26.750 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 6.455 1.760 9.870 1.885 ;
        RECT 12.970 1.760 18.650 1.885 ;
        RECT -0.430 -0.430 26.750 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 1.140 ;
        RECT 5.550 0.300 5.780 1.025 ;
        RECT 7.865 0.300 8.095 1.045 ;
        RECT 13.120 0.300 13.480 0.915 ;
        RECT 21.475 0.300 21.705 0.890 ;
        RECT 23.315 0.300 23.545 0.905 ;
        RECT 25.595 0.300 25.825 0.905 ;
        RECT 0.000 -0.300 26.320 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 6.085 3.160 7.360 3.390 ;
        RECT 0.245 2.615 0.475 3.040 ;
        RECT 3.270 2.745 4.120 2.975 ;
        RECT 3.890 2.655 4.120 2.745 ;
        RECT 6.085 2.655 6.315 3.160 ;
        RECT 7.130 3.120 7.360 3.160 ;
        RECT 8.205 3.160 9.835 3.390 ;
        RECT 11.265 3.215 12.780 3.390 ;
        RECT 13.760 3.215 15.230 3.390 ;
        RECT 11.265 3.160 15.230 3.215 ;
        RECT 8.205 3.120 8.435 3.160 ;
        RECT 7.130 2.890 8.435 3.120 ;
        RECT 0.245 2.385 2.855 2.615 ;
        RECT 3.890 2.420 6.315 2.655 ;
        RECT 6.610 2.620 6.840 2.890 ;
        RECT 6.610 2.385 8.535 2.620 ;
        RECT 0.245 0.780 0.475 2.385 ;
        RECT 2.625 1.535 2.855 2.385 ;
        RECT 4.630 1.535 4.860 1.740 ;
        RECT 2.625 1.305 4.860 1.535 ;
        RECT 5.090 1.260 6.240 1.490 ;
        RECT 6.945 1.275 7.175 2.385 ;
        RECT 8.305 1.910 8.535 2.385 ;
        RECT 8.885 2.035 9.115 2.890 ;
        RECT 9.605 2.485 9.835 3.160 ;
        RECT 12.550 2.985 13.990 3.160 ;
        RECT 10.800 2.295 11.030 2.870 ;
        RECT 10.800 2.065 14.255 2.295 ;
        RECT 14.485 2.220 14.715 2.930 ;
        RECT 15.000 2.680 15.230 3.160 ;
        RECT 16.050 3.115 17.250 3.345 ;
        RECT 16.050 2.680 16.280 3.115 ;
        RECT 15.000 2.450 16.280 2.680 ;
        RECT 16.510 2.220 16.740 2.885 ;
        RECT 8.885 1.800 10.390 2.035 ;
        RECT 5.090 1.075 5.320 1.260 ;
        RECT 3.250 0.845 5.320 1.075 ;
        RECT 6.010 0.760 6.240 1.260 ;
        RECT 6.835 0.990 7.175 1.275 ;
        RECT 7.405 1.295 8.680 1.530 ;
        RECT 7.405 0.760 7.635 1.295 ;
        RECT 6.010 0.530 7.635 0.760 ;
        RECT 8.450 0.760 8.680 1.295 ;
        RECT 9.150 0.990 9.490 1.800 ;
        RECT 9.925 0.760 10.155 0.980 ;
        RECT 8.450 0.530 10.155 0.760 ;
        RECT 11.045 0.620 11.275 2.065 ;
        RECT 14.485 1.990 16.740 2.220 ;
        RECT 17.020 2.065 17.250 3.115 ;
        RECT 17.530 3.115 19.240 3.345 ;
        RECT 14.485 1.835 14.715 1.990 ;
        RECT 11.625 1.375 11.855 1.700 ;
        RECT 12.475 1.605 14.715 1.835 ;
        RECT 11.625 1.145 14.330 1.375 ;
        RECT 14.100 0.760 14.330 1.145 ;
        RECT 15.470 0.990 15.810 1.990 ;
        RECT 17.530 1.760 17.760 3.115 ;
        RECT 18.550 2.315 18.780 2.885 ;
        RECT 19.010 2.735 19.240 3.115 ;
        RECT 20.055 3.160 21.330 3.390 ;
        RECT 20.055 2.735 20.285 3.160 ;
        RECT 19.010 2.505 20.285 2.735 ;
        RECT 16.090 0.760 16.320 1.740 ;
        RECT 16.590 1.525 17.760 1.760 ;
        RECT 17.990 2.275 18.780 2.315 ;
        RECT 17.990 2.045 19.280 2.275 ;
        RECT 16.590 0.990 16.930 1.525 ;
        RECT 17.990 1.265 18.220 2.045 ;
        RECT 17.710 0.990 18.220 1.265 ;
        RECT 18.450 0.760 18.820 1.815 ;
        RECT 14.100 0.530 18.820 0.760 ;
        RECT 19.050 0.760 19.280 2.045 ;
        RECT 20.525 0.760 20.865 2.930 ;
        RECT 21.100 2.735 21.330 3.160 ;
        RECT 21.100 2.505 22.540 2.735 ;
        RECT 21.115 1.725 21.345 2.170 ;
        RECT 22.200 1.960 22.540 2.505 ;
        RECT 22.800 2.095 23.030 3.380 ;
        RECT 22.800 1.825 25.300 2.095 ;
        RECT 22.800 1.725 23.030 1.825 ;
        RECT 21.115 1.495 23.030 1.725 ;
        RECT 19.050 0.530 20.865 0.760 ;
        RECT 22.595 0.655 23.030 1.495 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffsnq_2
MACRO gf180mcu_fd_sc_mcu7t5v0__sdffsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffsnq_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 29.680 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.408000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.410 1.770 4.430 2.150 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.816000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 0.595 1.030 2.150 ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.080500 ;
    PORT
      LAYER Metal1 ;
        RECT 20.075 1.210 21.230 1.590 ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.408000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.825 0.595 2.150 2.150 ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.686500 ;
    PORT
      LAYER Metal1 ;
        RECT 6.210 1.770 7.790 2.150 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.305500 ;
    PORT
      LAYER Metal1 ;
        RECT 25.310 2.290 25.640 3.380 ;
        RECT 27.440 2.290 27.910 3.380 ;
        RECT 25.310 2.055 27.910 2.290 ;
        RECT 27.440 1.345 27.910 2.055 ;
        RECT 25.310 1.115 27.910 1.345 ;
        RECT 25.310 0.805 25.540 1.115 ;
        RECT 27.440 0.595 27.910 1.115 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 29.680 4.220 ;
        RECT 1.260 2.845 1.600 3.620 ;
        RECT 5.250 3.305 5.590 3.620 ;
        RECT 8.100 3.350 8.440 3.620 ;
        RECT 13.510 3.360 13.850 3.620 ;
        RECT 15.985 2.930 16.215 3.620 ;
        RECT 19.930 2.660 20.270 3.620 ;
        RECT 22.285 2.530 22.515 3.620 ;
        RECT 24.325 2.530 24.555 3.620 ;
        RECT 26.380 2.530 26.610 3.620 ;
        RECT 28.570 2.530 28.800 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 30.110 4.350 ;
        RECT -0.430 1.760 5.965 1.885 ;
        RECT 21.345 1.760 30.110 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 5.965 1.760 21.345 1.885 ;
        RECT -0.430 -0.430 30.110 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.300 1.595 1.160 ;
        RECT 5.450 0.300 5.790 0.475 ;
        RECT 8.070 0.300 8.410 0.475 ;
        RECT 13.850 0.300 14.190 0.915 ;
        RECT 21.950 0.300 22.180 1.020 ;
        RECT 24.190 0.300 24.420 1.145 ;
        RECT 26.375 0.300 26.715 0.750 ;
        RECT 28.670 0.300 28.900 1.145 ;
        RECT 0.000 -0.300 29.680 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 5.820 3.160 7.790 3.390 ;
        RECT 0.245 2.615 0.475 3.140 ;
        RECT 5.820 3.075 6.050 3.160 ;
        RECT 3.270 2.845 6.050 3.075 ;
        RECT 7.560 3.120 7.790 3.160 ;
        RECT 8.865 3.120 10.850 3.295 ;
        RECT 7.560 3.065 10.850 3.120 ;
        RECT 7.560 2.890 9.095 3.065 ;
        RECT 6.785 2.660 7.070 2.835 ;
        RECT 0.245 2.385 5.065 2.615 ;
        RECT 6.785 2.430 9.045 2.660 ;
        RECT 9.395 2.495 9.995 2.835 ;
        RECT 10.510 2.655 10.850 3.065 ;
        RECT 12.110 3.130 12.450 3.355 ;
        RECT 14.320 3.160 15.710 3.390 ;
        RECT 14.320 3.130 14.550 3.160 ;
        RECT 0.245 0.780 0.475 2.385 ;
        RECT 2.600 2.105 2.830 2.385 ;
        RECT 4.725 1.455 5.065 2.385 ;
        RECT 8.815 1.395 9.045 2.430 ;
        RECT 6.510 1.165 9.045 1.395 ;
        RECT 9.710 2.280 9.995 2.495 ;
        RECT 9.710 2.045 11.290 2.280 ;
        RECT 3.270 0.935 3.610 1.095 ;
        RECT 6.510 0.990 6.850 1.165 ;
        RECT 9.710 0.990 10.050 2.045 ;
        RECT 11.585 1.960 11.815 3.015 ;
        RECT 12.110 2.900 14.550 3.130 ;
        RECT 14.910 2.425 15.250 2.780 ;
        RECT 15.480 2.700 15.710 3.160 ;
        RECT 16.700 3.040 17.990 3.310 ;
        RECT 16.700 2.700 16.930 3.040 ;
        RECT 15.480 2.465 16.930 2.700 ;
        RECT 12.850 2.190 15.250 2.425 ;
        RECT 14.965 2.040 15.250 2.190 ;
        RECT 17.170 2.040 17.510 2.810 ;
        RECT 18.245 2.105 18.475 2.890 ;
        RECT 11.585 1.725 14.670 1.960 ;
        RECT 14.965 1.805 17.510 2.040 ;
        RECT 17.810 1.875 18.475 2.105 ;
        RECT 19.265 2.430 19.495 2.890 ;
        RECT 21.005 2.430 21.235 2.835 ;
        RECT 19.265 2.200 21.235 2.430 ;
        RECT 3.270 0.760 6.250 0.935 ;
        RECT 7.610 0.760 9.315 0.935 ;
        RECT 10.665 0.760 10.895 0.970 ;
        RECT 3.270 0.705 10.895 0.760 ;
        RECT 6.020 0.530 7.840 0.705 ;
        RECT 9.085 0.530 10.895 0.705 ;
        RECT 11.785 0.680 12.015 1.725 ;
        RECT 12.310 1.260 14.975 1.495 ;
        RECT 14.745 0.760 14.975 1.260 ;
        RECT 16.030 0.990 16.370 1.805 ;
        RECT 17.810 1.220 18.040 1.875 ;
        RECT 19.265 1.220 19.495 2.200 ;
        RECT 23.305 2.195 23.535 3.380 ;
        RECT 21.530 1.965 23.535 2.195 ;
        RECT 23.070 1.805 23.535 1.965 ;
        RECT 21.490 1.450 22.775 1.685 ;
        RECT 23.070 1.575 27.105 1.805 ;
        RECT 17.150 0.990 18.040 1.220 ;
        RECT 18.270 0.990 19.770 1.220 ;
        RECT 17.810 0.760 18.040 0.990 ;
        RECT 21.490 0.760 21.720 1.450 ;
        RECT 23.070 0.805 23.300 1.575 ;
        RECT 14.745 0.530 16.810 0.760 ;
        RECT 17.810 0.530 21.720 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffsnq_4
MACRO gf180mcu_fd_sc_mcu7t5v0__tieh
  CLASS core TIEHIGH ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__tieh ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.220 2.305 1.580 3.390 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 2.240 4.220 ;
        RECT 0.250 2.360 0.480 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 2.670 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 0.300 0.480 1.160 ;
        RECT 0.000 -0.300 2.240 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.875 1.335 1.600 1.570 ;
        RECT 1.370 0.530 1.600 1.335 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__tieh
MACRO gf180mcu_fd_sc_mcu7t5v0__tiel
  CLASS core TIELOW ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__tiel ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.220 0.530 1.595 1.650 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 2.240 4.220 ;
        RECT 0.345 2.345 0.575 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 2.670 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 1.160 ;
        RECT 0.000 -0.300 2.240 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.365 2.185 1.595 3.390 ;
        RECT 0.870 1.950 1.595 2.185 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__tiel
MACRO gf180mcu_fd_sc_mcu7t5v0__xnor2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xnor2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.535500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.815 1.825 4.570 2.095 ;
        RECT 1.815 1.450 2.220 1.825 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.535500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.305 2.385 5.455 2.655 ;
        RECT 1.305 1.855 1.535 2.385 ;
        RECT 0.910 1.625 1.535 1.855 ;
        RECT 5.185 1.740 5.455 2.385 ;
        RECT 5.185 1.510 6.010 1.740 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.456350 ;
    PORT
      LAYER Metal1 ;
        RECT 3.305 2.945 6.020 3.215 ;
        RECT 5.745 2.215 6.020 2.945 ;
        RECT 5.745 1.980 6.580 2.215 ;
        RECT 6.290 1.220 6.580 1.980 ;
        RECT 4.980 0.990 6.580 1.220 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.280 4.220 ;
        RECT 0.385 2.720 0.615 3.620 ;
        RECT 2.650 2.930 2.990 3.620 ;
        RECT 6.305 2.690 6.535 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 7.710 4.350 ;
        RECT -0.430 1.760 4.630 1.885 ;
        RECT 5.730 1.760 7.710 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 4.630 1.760 5.730 1.885 ;
        RECT -0.430 -0.430 7.710 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.370 0.300 2.710 0.760 ;
        RECT 0.000 -0.300 7.280 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.845 2.945 1.780 3.215 ;
        RECT 0.845 2.415 1.075 2.945 ;
        RECT 0.330 2.180 1.075 2.415 ;
        RECT 0.330 1.220 0.615 2.180 ;
        RECT 3.105 1.220 3.445 1.565 ;
        RECT 0.330 0.990 3.445 1.220 ;
        RECT 0.330 0.530 0.670 0.990 ;
        RECT 3.630 0.530 6.690 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xnor2_1
MACRO gf180mcu_fd_sc_mcu7t5v0__xnor2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xnor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.600500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.825 1.825 4.105 2.095 ;
        RECT 1.825 1.570 2.290 1.825 ;
        RECT 3.855 1.745 4.105 1.825 ;
        RECT 3.855 1.255 4.480 1.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.600500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.260 2.470 4.520 2.660 ;
        RECT 1.260 2.325 5.475 2.470 ;
        RECT 1.260 1.885 1.535 2.325 ;
        RECT 4.290 2.235 5.475 2.325 ;
        RECT 0.835 1.655 1.535 1.885 ;
        RECT 5.215 1.785 5.475 2.235 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal1 ;
        RECT 7.585 0.600 8.265 3.380 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 9.520 4.220 ;
        RECT 2.435 2.915 2.665 3.620 ;
        RECT 6.545 2.530 6.775 3.620 ;
        RECT 8.685 2.530 8.915 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 9.950 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.300 0.475 0.825 ;
        RECT 2.485 0.300 2.715 0.825 ;
        RECT 5.825 0.300 6.055 0.915 ;
        RECT 6.545 0.300 6.775 0.915 ;
        RECT 8.785 0.300 9.015 1.115 ;
        RECT 0.000 -0.300 9.520 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 1.290 0.575 3.360 ;
        RECT 3.640 3.160 6.110 3.390 ;
        RECT 4.750 2.700 5.935 2.930 ;
        RECT 3.040 1.365 3.535 1.595 ;
        RECT 5.705 1.555 5.935 2.700 ;
        RECT 6.920 1.555 7.290 2.110 ;
        RECT 3.040 1.290 3.270 1.365 ;
        RECT 0.345 1.055 3.270 1.290 ;
        RECT 4.810 1.155 7.290 1.555 ;
        RECT 1.310 0.530 1.650 1.055 ;
        RECT 4.810 0.820 5.040 1.155 ;
        RECT 3.640 0.590 5.040 0.820 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xnor2_2
MACRO gf180mcu_fd_sc_mcu7t5v0__xnor2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xnor2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.760 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.498000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.830 2.010 4.060 2.120 ;
        RECT 1.830 1.795 4.550 2.010 ;
        RECT 1.830 1.580 2.225 1.795 ;
        RECT 3.785 1.660 4.550 1.795 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.498000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.260 2.470 4.520 2.680 ;
        RECT 1.260 2.360 5.070 2.470 ;
        RECT 1.260 2.095 1.535 2.360 ;
        RECT 4.290 2.240 5.070 2.360 ;
        RECT 0.755 1.810 1.535 2.095 ;
        RECT 4.840 2.100 5.070 2.240 ;
        RECT 4.840 1.810 5.630 2.100 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.243600 ;
    PORT
      LAYER Metal1 ;
        RECT 7.610 2.700 7.950 3.380 ;
        RECT 9.800 2.700 10.140 3.380 ;
        RECT 7.610 2.360 11.060 2.700 ;
        RECT 10.775 1.430 11.060 2.360 ;
        RECT 7.665 1.195 11.060 1.430 ;
        RECT 7.665 0.530 7.895 1.195 ;
        RECT 9.905 0.530 10.135 1.195 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 11.760 4.220 ;
        RECT 2.665 2.940 2.895 3.620 ;
        RECT 6.645 2.530 6.875 3.620 ;
        RECT 8.735 3.015 8.965 3.620 ;
        RECT 10.925 3.015 11.155 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 12.190 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.190 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 0.760 ;
        RECT 2.430 0.300 2.770 0.760 ;
        RECT 5.825 0.300 6.055 0.915 ;
        RECT 6.545 0.300 6.775 0.915 ;
        RECT 8.785 0.300 9.015 0.915 ;
        RECT 11.025 0.300 11.255 0.915 ;
        RECT 0.000 -0.300 11.760 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.575 3.160 6.110 3.390 ;
        RECT 0.230 1.225 0.525 2.720 ;
        RECT 4.750 2.700 6.240 2.930 ;
        RECT 6.010 1.895 6.240 2.700 ;
        RECT 6.010 1.665 10.500 1.895 ;
        RECT 3.000 1.225 3.400 1.555 ;
        RECT 6.010 1.430 6.240 1.665 ;
        RECT 0.230 0.990 3.400 1.225 ;
        RECT 3.785 1.195 6.240 1.430 ;
        RECT 1.310 0.530 1.650 0.990 ;
        RECT 3.785 0.530 4.015 1.195 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xnor2_4
MACRO gf180mcu_fd_sc_mcu7t5v0__xnor3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xnor3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.440 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.892000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.770 1.825 3.900 2.095 ;
        RECT 1.770 1.455 2.225 1.825 ;
        RECT 3.670 1.690 3.900 1.825 ;
        RECT 3.670 1.455 4.770 1.690 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.892000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.870 2.385 4.360 2.655 ;
        RECT 4.130 2.150 4.360 2.385 ;
        RECT 4.130 1.920 5.620 2.150 ;
        RECT 5.175 1.595 5.620 1.920 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.535500 ;
    PORT
      LAYER Metal1 ;
        RECT 8.085 1.825 10.765 2.095 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.511100 ;
    PORT
      LAYER Metal1 ;
        RECT 9.570 2.920 12.215 3.240 ;
        RECT 11.880 2.680 12.215 2.920 ;
        RECT 11.880 2.360 12.760 2.680 ;
        RECT 12.440 1.580 12.760 2.360 ;
        RECT 11.170 0.990 12.760 1.580 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 13.440 4.220 ;
        RECT 2.370 2.900 2.730 3.620 ;
        RECT 6.545 2.840 6.775 3.620 ;
        RECT 8.760 2.815 9.100 3.620 ;
        RECT 12.465 3.015 12.695 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 13.870 4.350 ;
        RECT -0.430 1.760 10.790 1.885 ;
        RECT 11.890 1.760 13.870 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 10.790 1.760 11.890 1.885 ;
        RECT -0.430 -0.430 13.870 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 0.760 ;
        RECT 2.430 0.300 2.770 0.760 ;
        RECT 5.770 0.300 6.110 0.760 ;
        RECT 8.530 0.300 8.870 0.760 ;
        RECT 0.000 -0.300 13.440 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 1.220 0.575 3.195 ;
        RECT 3.720 3.160 6.120 3.390 ;
        RECT 3.720 2.900 4.080 3.160 ;
        RECT 4.740 2.610 5.100 2.930 ;
        RECT 5.760 2.900 6.120 3.160 ;
        RECT 7.030 3.160 8.500 3.390 ;
        RECT 7.030 2.610 7.260 3.160 ;
        RECT 4.740 2.380 7.260 2.610 ;
        RECT 5.880 1.225 6.110 2.380 ;
        RECT 7.030 1.535 7.260 2.380 ;
        RECT 7.510 1.225 7.850 2.930 ;
        RECT 8.270 2.565 8.500 3.160 ;
        RECT 8.270 2.330 11.450 2.565 ;
        RECT 11.220 2.095 11.450 2.330 ;
        RECT 11.220 1.860 12.170 2.095 ;
        RECT 9.200 1.225 9.540 1.565 ;
        RECT 0.345 0.990 3.495 1.220 ;
        RECT 3.730 0.990 6.110 1.225 ;
        RECT 6.490 0.990 9.540 1.225 ;
        RECT 1.305 0.530 1.650 0.990 ;
        RECT 3.730 0.530 4.070 0.990 ;
        RECT 6.490 0.530 6.830 0.990 ;
        RECT 9.740 0.530 12.860 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xnor3_1
MACRO gf180mcu_fd_sc_mcu7t5v0__xnor3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xnor3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.680 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.904500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.935 1.265 4.905 1.535 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.904500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.825 2.385 4.240 2.655 ;
        RECT 3.935 2.100 4.240 2.385 ;
        RECT 3.935 1.815 5.715 2.100 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.598000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.300 1.815 10.425 2.095 ;
        RECT 10.170 1.610 10.425 1.815 ;
        RECT 10.170 1.210 11.075 1.610 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.795200 ;
    PORT
      LAYER Metal1 ;
        RECT 13.015 2.680 13.295 3.390 ;
        RECT 15.155 2.680 15.535 3.390 ;
        RECT 13.015 2.360 15.535 2.680 ;
        RECT 15.155 1.560 15.535 2.360 ;
        RECT 12.965 1.240 15.535 1.560 ;
        RECT 12.965 0.600 13.310 1.240 ;
        RECT 15.155 0.600 15.535 1.240 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 15.680 4.220 ;
        RECT 2.420 2.895 2.780 3.620 ;
        RECT 9.090 2.785 9.430 3.620 ;
        RECT 14.035 2.950 14.265 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 16.110 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 16.110 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 0.760 ;
        RECT 2.515 0.300 2.855 0.760 ;
        RECT 5.770 0.300 6.110 0.760 ;
        RECT 6.570 0.300 6.910 0.760 ;
        RECT 9.045 0.300 9.275 0.890 ;
        RECT 12.150 0.300 12.490 0.635 ;
        RECT 14.085 0.300 14.315 0.975 ;
        RECT 0.000 -0.300 15.680 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.345 1.225 0.575 3.190 ;
        RECT 3.720 3.155 6.055 3.390 ;
        RECT 3.720 2.895 4.080 3.155 ;
        RECT 4.750 2.565 5.090 2.925 ;
        RECT 5.760 2.840 6.055 3.155 ;
        RECT 6.285 3.155 8.065 3.390 ;
        RECT 10.045 3.160 12.575 3.390 ;
        RECT 6.285 2.565 6.515 3.155 ;
        RECT 4.750 2.335 6.515 2.565 ;
        RECT 1.365 1.765 3.570 1.995 ;
        RECT 1.365 1.225 1.650 1.765 ;
        RECT 0.345 0.990 1.650 1.225 ;
        RECT 6.285 1.225 6.515 2.335 ;
        RECT 6.745 2.095 7.085 2.925 ;
        RECT 7.835 2.555 8.065 3.155 ;
        RECT 11.115 2.700 12.575 2.930 ;
        RECT 7.835 2.470 10.885 2.555 ;
        RECT 7.835 2.325 11.995 2.470 ;
        RECT 10.655 2.240 11.995 2.325 ;
        RECT 6.745 1.860 8.030 2.095 ;
        RECT 7.690 1.380 8.030 1.860 ;
        RECT 11.765 1.715 11.995 2.240 ;
        RECT 12.345 2.045 12.575 2.700 ;
        RECT 12.345 1.815 14.915 2.045 ;
        RECT 9.515 1.380 9.905 1.555 ;
        RECT 6.285 1.220 7.435 1.225 ;
        RECT 1.310 0.530 1.650 0.990 ;
        RECT 5.230 0.990 7.435 1.220 ;
        RECT 7.690 1.150 9.905 1.380 ;
        RECT 5.230 0.760 5.460 0.990 ;
        RECT 3.730 0.530 5.460 0.760 ;
        RECT 7.690 0.530 8.030 1.150 ;
        RECT 12.345 1.095 12.575 1.815 ;
        RECT 11.405 0.865 12.575 1.095 ;
        RECT 11.405 0.765 11.710 0.865 ;
        RECT 10.035 0.530 11.710 0.765 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xnor3_2
MACRO gf180mcu_fd_sc_mcu7t5v0__xnor3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xnor3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.920 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.804500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.880 1.240 4.420 1.535 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.804500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.875 2.265 3.890 2.495 ;
        RECT 0.875 1.565 1.105 2.265 ;
        RECT 3.450 2.095 3.890 2.265 ;
        RECT 3.450 1.820 5.260 2.095 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.510500 ;
    PORT
      LAYER Metal1 ;
        RECT 8.175 1.800 10.275 2.095 ;
        RECT 10.020 1.565 10.275 1.800 ;
        RECT 10.020 1.255 11.150 1.565 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.978000 ;
    PORT
      LAYER Metal1 ;
        RECT 12.940 2.680 13.170 3.380 ;
        RECT 15.030 2.680 15.260 3.380 ;
        RECT 17.220 2.680 17.775 3.380 ;
        RECT 12.940 2.360 17.775 2.680 ;
        RECT 17.320 1.535 17.775 2.360 ;
        RECT 12.840 1.260 17.775 1.535 ;
        RECT 12.840 0.655 13.070 1.260 ;
        RECT 15.080 0.655 15.310 1.260 ;
        RECT 17.320 0.600 17.775 1.260 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 17.920 4.220 ;
        RECT 2.330 2.725 2.670 3.620 ;
        RECT 8.965 2.785 9.305 3.620 ;
        RECT 13.960 3.015 14.190 3.620 ;
        RECT 16.150 3.015 16.380 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 18.350 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 18.350 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 0.760 ;
        RECT 2.430 0.300 2.770 0.760 ;
        RECT 5.590 0.300 6.740 0.760 ;
        RECT 8.915 0.300 9.145 0.840 ;
        RECT 12.025 0.300 12.365 0.640 ;
        RECT 13.960 0.300 14.190 0.905 ;
        RECT 16.200 0.300 16.430 0.905 ;
        RECT 0.000 -0.300 17.920 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.550 3.160 6.165 3.390 ;
        RECT 0.345 1.225 0.575 3.015 ;
        RECT 3.550 2.725 3.890 3.160 ;
        RECT 4.570 2.555 4.910 2.930 ;
        RECT 5.825 2.725 6.165 3.160 ;
        RECT 6.395 3.160 8.390 3.390 ;
        RECT 9.895 3.160 12.375 3.390 ;
        RECT 4.570 2.495 5.670 2.555 ;
        RECT 6.395 2.495 6.625 3.160 ;
        RECT 4.570 2.325 6.625 2.495 ;
        RECT 5.440 2.265 6.625 2.325 ;
        RECT 1.420 1.765 3.220 2.035 ;
        RECT 1.420 1.225 1.650 1.765 ;
        RECT 6.395 1.535 6.625 2.265 ;
        RECT 6.905 2.095 7.245 2.930 ;
        RECT 8.115 2.555 8.390 3.160 ;
        RECT 10.915 2.700 12.375 2.930 ;
        RECT 8.115 2.325 10.735 2.555 ;
        RECT 10.505 2.180 10.735 2.325 ;
        RECT 6.905 1.800 7.860 2.095 ;
        RECT 10.505 1.820 11.760 2.180 ;
        RECT 12.145 1.995 12.375 2.700 ;
        RECT 0.345 0.990 1.650 1.225 ;
        RECT 1.310 0.530 1.650 0.990 ;
        RECT 5.115 1.300 7.275 1.535 ;
        RECT 7.520 1.305 7.860 1.800 ;
        RECT 12.145 1.765 17.060 1.995 ;
        RECT 9.405 1.305 9.745 1.560 ;
        RECT 12.145 1.485 12.375 1.765 ;
        RECT 5.115 0.760 5.345 1.300 ;
        RECT 3.550 0.530 5.345 0.760 ;
        RECT 7.520 1.075 9.745 1.305 ;
        RECT 11.565 1.255 12.375 1.485 ;
        RECT 7.520 0.530 7.860 1.075 ;
        RECT 11.565 0.760 11.795 1.255 ;
        RECT 9.895 0.530 11.795 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xnor3_4
MACRO gf180mcu_fd_sc_mcu7t5v0__xor2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xor2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.598000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.875 1.820 4.015 2.100 ;
        RECT 3.785 1.570 4.015 1.820 ;
        RECT 3.785 1.340 4.525 1.570 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.598000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.880 2.560 2.325 2.730 ;
        RECT 0.880 2.330 4.495 2.560 ;
        RECT 0.880 1.690 1.560 2.330 ;
        RECT 4.255 2.155 4.495 2.330 ;
        RECT 4.255 1.800 5.490 2.155 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.060800 ;
    PORT
      LAYER Metal1 ;
        RECT 4.750 2.695 6.040 2.925 ;
        RECT 5.720 1.110 6.040 2.695 ;
        RECT 3.785 0.875 6.040 1.110 ;
        RECT 3.785 0.530 4.015 0.875 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 6.720 4.220 ;
        RECT 2.710 2.790 3.050 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 7.150 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.150 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 0.760 ;
        RECT 2.610 0.300 2.950 0.760 ;
        RECT 5.770 0.300 6.110 0.635 ;
        RECT 0.000 -0.300 6.720 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.290 1.290 0.630 3.350 ;
        RECT 3.590 3.155 6.120 3.390 ;
        RECT 3.170 1.290 3.510 1.555 ;
        RECT 0.290 0.990 3.510 1.290 ;
        RECT 1.310 0.530 1.650 0.990 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xor2_1
MACRO gf180mcu_fd_sc_mcu7t5v0__xor2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.535500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.595 1.795 4.565 2.095 ;
        RECT 2.595 1.680 2.870 1.795 ;
        RECT 1.850 1.450 2.870 1.680 ;
        RECT 4.270 1.265 4.565 1.795 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.535500 ;
    PORT
      LAYER Metal1 ;
        RECT 3.375 2.555 5.105 2.680 ;
        RECT 2.035 2.325 5.105 2.555 ;
        RECT 2.035 2.140 2.315 2.325 ;
        RECT 0.915 1.910 2.315 2.140 ;
        RECT 4.830 2.120 5.105 2.325 ;
        RECT 0.915 1.800 1.610 1.910 ;
        RECT 4.830 1.800 6.225 2.120 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.060800 ;
    PORT
      LAYER Metal1 ;
        RECT 8.195 2.680 8.560 3.380 ;
        RECT 8.195 2.360 9.600 2.680 ;
        RECT 9.315 1.560 9.600 2.360 ;
        RECT 8.195 1.240 9.600 1.560 ;
        RECT 8.195 0.610 8.545 1.240 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 10.080 4.220 ;
        RECT 0.455 2.830 0.685 3.620 ;
        RECT 2.720 2.790 3.060 3.620 ;
        RECT 6.320 2.815 6.660 3.620 ;
        RECT 7.295 2.530 7.525 3.620 ;
        RECT 9.335 2.940 9.565 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 10.510 4.350 ;
        RECT -0.430 1.760 4.700 1.885 ;
        RECT 5.800 1.760 10.510 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 4.700 1.760 5.800 1.885 ;
        RECT -0.430 -0.430 10.510 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.620 0.300 2.960 0.760 ;
        RECT 7.195 0.300 7.425 0.990 ;
        RECT 9.435 0.300 9.665 0.990 ;
        RECT 0.000 -0.300 10.080 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 1.475 2.600 1.705 3.350 ;
        RECT 3.600 2.990 5.630 3.220 ;
        RECT 0.400 2.370 1.705 2.600 ;
        RECT 5.400 2.580 5.630 2.990 ;
        RECT 0.400 1.220 0.680 2.370 ;
        RECT 5.400 2.350 6.770 2.580 ;
        RECT 6.540 2.095 6.770 2.350 ;
        RECT 6.540 1.820 9.080 2.095 ;
        RECT 3.180 1.220 3.520 1.555 ;
        RECT 6.540 1.220 6.770 1.820 ;
        RECT 0.400 0.990 3.520 1.220 ;
        RECT 5.070 0.990 6.770 1.220 ;
        RECT 0.400 0.530 0.740 0.990 ;
        RECT 3.650 0.530 6.770 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xor2_2
MACRO gf180mcu_fd_sc_mcu7t5v0__xor2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xor2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.320 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.448000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.935 1.825 4.525 2.095 ;
        RECT 4.225 1.230 4.525 1.825 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.448000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.000 2.555 5.025 2.680 ;
        RECT 1.425 2.325 5.025 2.555 ;
        RECT 1.425 2.100 1.700 2.325 ;
        RECT 0.860 1.810 1.700 2.100 ;
        RECT 4.795 2.120 5.025 2.325 ;
        RECT 4.795 1.800 6.180 2.120 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.243600 ;
    PORT
      LAYER Metal1 ;
        RECT 8.270 2.680 8.500 3.380 ;
        RECT 10.460 2.680 10.690 3.380 ;
        RECT 8.270 2.360 11.780 2.680 ;
        RECT 11.510 1.560 11.780 2.360 ;
        RECT 8.270 1.240 11.780 1.560 ;
        RECT 8.270 0.655 8.500 1.240 ;
        RECT 10.510 0.655 10.740 1.240 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 12.320 4.220 ;
        RECT 0.355 2.795 0.695 3.620 ;
        RECT 2.395 2.785 2.735 3.620 ;
        RECT 6.275 2.815 6.615 3.620 ;
        RECT 7.250 2.530 7.480 3.620 ;
        RECT 9.340 3.000 9.570 3.620 ;
        RECT 11.530 3.000 11.760 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 12.750 4.350 ;
        RECT -0.430 1.760 4.655 1.885 ;
        RECT 5.755 1.760 12.750 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 4.655 1.760 5.755 1.885 ;
        RECT -0.430 -0.430 12.750 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.575 0.300 2.915 0.760 ;
        RECT 7.150 0.300 7.380 0.905 ;
        RECT 9.390 0.300 9.620 0.985 ;
        RECT 11.630 0.300 11.860 0.985 ;
        RECT 0.000 -0.300 12.320 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.930 2.785 1.805 3.015 ;
        RECT 3.660 2.965 5.680 3.195 ;
        RECT 0.930 2.565 1.190 2.785 ;
        RECT 0.355 2.330 1.190 2.565 ;
        RECT 5.450 2.585 5.680 2.965 ;
        RECT 5.450 2.350 6.725 2.585 ;
        RECT 0.355 1.220 0.585 2.330 ;
        RECT 6.495 2.105 6.725 2.350 ;
        RECT 6.495 1.815 11.275 2.105 ;
        RECT 3.170 1.220 3.510 1.555 ;
        RECT 6.495 1.220 6.725 1.815 ;
        RECT 0.355 0.990 3.510 1.220 ;
        RECT 4.920 0.990 6.725 1.220 ;
        RECT 0.355 0.530 0.695 0.990 ;
        RECT 3.605 0.530 6.725 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xor2_4
MACRO gf180mcu_fd_sc_mcu7t5v0__xor3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xor3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.880 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.894500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.890 1.265 4.600 1.535 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.894500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.865 2.455 2.100 2.710 ;
        RECT 0.865 2.225 4.195 2.455 ;
        RECT 0.865 1.570 1.095 2.225 ;
        RECT 3.915 2.095 4.195 2.225 ;
        RECT 3.915 1.820 5.600 2.095 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.600500 ;
    PORT
      LAYER Metal1 ;
        RECT 8.205 1.825 10.205 2.100 ;
        RECT 8.205 1.455 8.545 1.825 ;
        RECT 9.975 1.560 10.205 1.825 ;
        RECT 9.975 1.265 11.110 1.560 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.060800 ;
    PORT
      LAYER Metal1 ;
        RECT 10.770 2.700 12.200 2.930 ;
        RECT 11.880 1.295 12.200 2.700 ;
        RECT 11.560 1.015 12.200 1.295 ;
        RECT 11.560 1.000 11.830 1.015 ;
        RECT 10.045 0.670 11.830 1.000 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 12.880 4.220 ;
        RECT 2.330 2.685 2.670 3.620 ;
        RECT 8.750 2.790 9.090 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.760 13.310 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 13.310 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 0.760 ;
        RECT 2.430 0.300 2.770 0.760 ;
        RECT 5.770 0.300 6.850 0.760 ;
        RECT 8.915 0.300 9.275 0.760 ;
        RECT 12.085 0.300 12.425 0.635 ;
        RECT 0.000 -0.300 12.880 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.730 3.160 6.055 3.390 ;
        RECT 0.345 1.305 0.575 2.980 ;
        RECT 3.730 2.755 4.070 3.160 ;
        RECT 4.750 2.555 5.090 2.915 ;
        RECT 5.825 2.815 6.055 3.160 ;
        RECT 6.285 3.160 7.925 3.390 ;
        RECT 9.640 3.160 12.160 3.390 ;
        RECT 6.285 2.555 6.515 3.160 ;
        RECT 4.750 2.325 6.515 2.555 ;
        RECT 1.385 1.765 3.510 1.995 ;
        RECT 1.385 1.305 1.650 1.765 ;
        RECT 5.880 1.305 6.110 2.325 ;
        RECT 6.745 1.765 6.975 2.925 ;
        RECT 7.695 2.560 7.925 3.160 ;
        RECT 7.695 2.470 10.585 2.560 ;
        RECT 7.695 2.330 11.585 2.470 ;
        RECT 10.395 2.240 11.585 2.330 ;
        RECT 6.745 1.535 7.930 1.765 ;
        RECT 11.350 1.760 11.585 2.240 ;
        RECT 0.345 1.070 1.650 1.305 ;
        RECT 1.310 0.530 1.650 1.070 ;
        RECT 5.195 1.070 7.390 1.305 ;
        RECT 7.625 1.220 7.930 1.535 ;
        RECT 9.395 1.220 9.745 1.555 ;
        RECT 5.195 0.760 5.425 1.070 ;
        RECT 3.700 0.530 5.425 0.760 ;
        RECT 7.625 0.990 9.745 1.220 ;
        RECT 7.625 0.530 7.965 0.990 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xor3_1
MACRO gf180mcu_fd_sc_mcu7t5v0__xor3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xor3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.240 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.892000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.050 1.265 4.535 1.535 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.892000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.075 2.455 2.275 2.660 ;
        RECT 1.075 2.225 4.065 2.455 ;
        RECT 1.075 1.490 1.305 2.225 ;
        RECT 3.835 2.095 4.065 2.225 ;
        RECT 3.835 1.765 5.095 2.095 ;
        RECT 4.800 1.720 5.095 1.765 ;
        RECT 4.800 1.485 5.695 1.720 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.535500 ;
    PORT
      LAYER Metal1 ;
        RECT 8.115 1.825 10.710 2.095 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.795200 ;
    PORT
      LAYER Metal1 ;
        RECT 13.290 2.680 13.520 3.360 ;
        RECT 15.240 2.680 15.760 3.360 ;
        RECT 13.290 2.360 15.760 2.680 ;
        RECT 15.460 1.560 15.760 2.360 ;
        RECT 13.290 1.240 15.760 1.560 ;
        RECT 13.290 0.655 13.520 1.240 ;
        RECT 15.530 0.655 15.760 1.240 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 16.240 4.220 ;
        RECT 2.725 2.735 3.065 3.620 ;
        RECT 6.525 2.680 6.810 3.620 ;
        RECT 8.775 2.795 9.135 3.620 ;
        RECT 11.990 3.280 12.355 3.620 ;
        RECT 14.310 3.015 14.540 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 16.670 4.350 ;
        RECT -0.430 1.760 10.795 1.885 ;
        RECT 11.895 1.760 16.670 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 10.795 1.760 11.895 1.885 ;
        RECT -0.430 -0.430 16.670 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.355 0.300 0.695 0.760 ;
        RECT 2.595 0.300 2.935 0.775 ;
        RECT 5.755 0.300 6.095 0.760 ;
        RECT 8.535 0.300 8.880 0.760 ;
        RECT 14.410 0.300 14.640 0.905 ;
        RECT 0.000 -0.300 16.240 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.735 3.160 6.070 3.390 ;
        RECT 0.510 1.220 0.740 3.030 ;
        RECT 3.735 2.735 4.095 3.160 ;
        RECT 4.720 2.605 5.555 2.835 ;
        RECT 5.785 2.680 6.070 3.160 ;
        RECT 7.040 3.010 8.445 3.240 ;
        RECT 5.325 2.220 5.555 2.605 ;
        RECT 7.040 2.220 7.270 3.010 ;
        RECT 1.535 1.765 3.560 1.995 ;
        RECT 5.325 1.990 7.270 2.220 ;
        RECT 1.535 1.220 1.815 1.765 ;
        RECT 7.010 1.220 7.270 1.990 ;
        RECT 0.510 0.990 1.815 1.220 ;
        RECT 1.475 0.530 1.815 0.990 ;
        RECT 5.240 0.990 7.270 1.220 ;
        RECT 7.545 1.220 7.885 2.780 ;
        RECT 8.160 2.565 8.445 3.010 ;
        RECT 9.750 2.815 12.355 3.050 ;
        RECT 8.160 2.330 11.335 2.565 ;
        RECT 11.105 1.900 11.335 2.330 ;
        RECT 12.125 2.095 12.355 2.815 ;
        RECT 11.105 1.670 11.760 1.900 ;
        RECT 12.125 1.825 15.210 2.095 ;
        RECT 9.270 1.220 9.610 1.555 ;
        RECT 12.125 1.220 12.355 1.825 ;
        RECT 7.545 0.990 9.610 1.220 ;
        RECT 11.170 0.990 12.355 1.220 ;
        RECT 5.240 0.760 5.470 0.990 ;
        RECT 7.545 0.760 7.885 0.990 ;
        RECT 3.625 0.530 5.470 0.760 ;
        RECT 6.485 0.530 7.885 0.760 ;
        RECT 9.795 0.530 12.865 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xor3_2
MACRO gf180mcu_fd_sc_mcu7t5v0__xor3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xor3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.480 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.804500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.880 1.265 4.360 1.535 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.804500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.865 2.455 2.100 2.710 ;
        RECT 0.865 2.225 3.875 2.455 ;
        RECT 0.865 1.600 1.105 2.225 ;
        RECT 3.645 2.095 3.875 2.225 ;
        RECT 3.645 1.820 4.895 2.095 ;
        RECT 4.615 1.790 4.895 1.820 ;
        RECT 4.615 1.560 5.360 1.790 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.435500 ;
    PORT
      LAYER Metal1 ;
        RECT 7.910 1.820 10.600 2.115 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.978000 ;
    PORT
      LAYER Metal1 ;
        RECT 13.025 2.680 13.505 3.315 ;
        RECT 15.265 2.680 15.690 3.315 ;
        RECT 17.370 2.680 17.815 3.325 ;
        RECT 13.025 2.360 17.815 2.680 ;
        RECT 17.480 1.560 17.815 2.360 ;
        RECT 13.025 1.240 17.815 1.560 ;
        RECT 13.025 0.600 13.335 1.240 ;
        RECT 15.265 0.600 15.575 1.240 ;
        RECT 17.505 0.600 17.815 1.240 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 18.480 4.220 ;
        RECT 2.330 2.685 2.670 3.620 ;
        RECT 6.365 2.485 6.595 3.620 ;
        RECT 8.570 2.805 8.910 3.620 ;
        RECT 12.230 3.285 12.570 3.620 ;
        RECT 14.225 2.940 14.455 3.620 ;
        RECT 16.415 2.940 16.645 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.885 18.910 4.350 ;
        RECT -0.430 1.760 10.610 1.885 ;
        RECT 11.710 1.760 18.910 1.885 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 10.610 1.760 11.710 1.885 ;
        RECT -0.430 -0.430 18.910 1.760 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.190 0.300 0.530 0.760 ;
        RECT 2.430 0.300 2.770 0.760 ;
        RECT 5.590 0.300 5.930 0.760 ;
        RECT 8.350 0.300 8.690 0.775 ;
        RECT 14.225 0.300 14.455 0.850 ;
        RECT 16.465 0.300 16.695 0.840 ;
        RECT 0.000 -0.300 18.480 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 3.550 3.160 5.875 3.390 ;
        RECT 0.345 1.355 0.575 2.980 ;
        RECT 3.550 2.685 3.890 3.160 ;
        RECT 4.570 2.685 5.370 2.915 ;
        RECT 5.140 2.260 5.370 2.685 ;
        RECT 5.645 2.610 5.875 3.160 ;
        RECT 6.885 3.140 8.205 3.390 ;
        RECT 5.140 2.025 5.935 2.260 ;
        RECT 1.350 1.765 3.410 1.995 ;
        RECT 1.350 1.355 1.580 1.765 ;
        RECT 0.345 1.120 1.580 1.355 ;
        RECT 5.705 1.305 5.935 2.025 ;
        RECT 6.885 1.305 7.115 3.140 ;
        RECT 0.835 0.760 1.085 1.120 ;
        RECT 5.035 1.075 7.115 1.305 ;
        RECT 7.385 1.585 7.615 2.845 ;
        RECT 7.970 2.575 8.205 3.140 ;
        RECT 9.635 2.815 12.575 3.050 ;
        RECT 7.970 2.345 11.995 2.575 ;
        RECT 11.765 1.695 11.995 2.345 ;
        RECT 12.345 2.095 12.575 2.815 ;
        RECT 12.345 1.825 17.225 2.095 ;
        RECT 7.385 1.350 9.555 1.585 ;
        RECT 5.035 0.760 5.265 1.075 ;
        RECT 7.385 0.765 7.615 1.350 ;
        RECT 12.345 1.220 12.575 1.825 ;
        RECT 10.980 0.990 12.575 1.220 ;
        RECT 0.835 0.530 1.650 0.760 ;
        RECT 3.550 0.530 5.265 0.760 ;
        RECT 6.310 0.530 7.615 0.765 ;
        RECT 9.560 0.530 12.680 0.760 ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xor3_4
END LIBRARY