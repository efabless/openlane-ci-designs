module user_proj_example (wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    vdd,
    vss,
    io_in,
    io_oeb,
    io_out,
    irq,
    la_data_in,
    la_data_out,
    la_oenb,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input vdd;
 input vss;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [2:0] irq;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;


 gf180mcu_fd_sc_mcu9t5v0__tieh _000_ (.Z(wbs_ack_o),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _001_ (.ZN(io_oeb[10]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _002_ (.ZN(io_oeb[11]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _003_ (.ZN(io_oeb[12]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _004_ (.ZN(io_oeb[13]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _005_ (.ZN(io_oeb[14]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _006_ (.ZN(io_oeb[15]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _007_ (.ZN(io_oeb[16]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _008_ (.ZN(io_oeb[17]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _009_ (.ZN(io_oeb[18]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _010_ (.ZN(io_oeb[19]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _011_ (.ZN(io_oeb[20]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _012_ (.ZN(io_oeb[21]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _013_ (.ZN(io_oeb[22]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _014_ (.ZN(io_oeb[23]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _015_ (.ZN(io_oeb[24]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _016_ (.ZN(io_oeb[25]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _017_ (.ZN(io_oeb[26]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _018_ (.ZN(io_oeb[27]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _019_ (.ZN(io_oeb[28]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _020_ (.ZN(io_oeb[29]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _021_ (.ZN(io_oeb[30]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _022_ (.ZN(io_oeb[31]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _023_ (.ZN(io_oeb[32]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _024_ (.ZN(io_oeb[33]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _025_ (.ZN(io_oeb[34]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _026_ (.ZN(io_oeb[35]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _027_ (.ZN(io_oeb[36]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _028_ (.ZN(io_oeb[37]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _029_ (.ZN(io_out[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _030_ (.ZN(io_out[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _031_ (.ZN(io_out[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _032_ (.ZN(io_out[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _033_ (.ZN(io_out[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _034_ (.ZN(io_out[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _035_ (.ZN(io_out[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _036_ (.ZN(io_out[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _037_ (.ZN(io_out[8]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _038_ (.ZN(io_out[9]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _039_ (.ZN(io_out[10]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _040_ (.ZN(io_out[11]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _041_ (.ZN(io_out[12]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _042_ (.ZN(io_out[13]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _043_ (.ZN(io_out[14]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _044_ (.ZN(io_out[15]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _045_ (.ZN(io_out[16]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _046_ (.ZN(io_out[17]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _047_ (.ZN(io_out[18]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _048_ (.ZN(io_out[19]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _049_ (.ZN(io_out[20]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _050_ (.ZN(io_out[21]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _051_ (.ZN(io_out[22]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _052_ (.ZN(io_out[23]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _053_ (.ZN(io_out[24]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _054_ (.ZN(io_out[25]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _055_ (.ZN(io_out[26]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _056_ (.ZN(io_out[27]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _057_ (.ZN(io_out[28]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _058_ (.ZN(io_out[29]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _059_ (.ZN(io_out[30]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _060_ (.ZN(io_out[31]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _061_ (.ZN(io_out[32]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _062_ (.ZN(io_out[33]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _063_ (.ZN(io_out[34]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _064_ (.ZN(io_out[35]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _065_ (.ZN(io_out[36]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _066_ (.ZN(io_out[37]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _067_ (.ZN(irq[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _068_ (.ZN(irq[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _069_ (.ZN(irq[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _070_ (.ZN(la_data_out[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _071_ (.ZN(la_data_out[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _072_ (.ZN(la_data_out[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _073_ (.ZN(la_data_out[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _074_ (.ZN(la_data_out[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _075_ (.ZN(la_data_out[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _076_ (.ZN(la_data_out[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _077_ (.ZN(la_data_out[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _078_ (.ZN(la_data_out[8]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _079_ (.ZN(la_data_out[9]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _080_ (.ZN(la_data_out[10]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _081_ (.ZN(la_data_out[11]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _082_ (.ZN(la_data_out[12]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _083_ (.ZN(la_data_out[13]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _084_ (.ZN(la_data_out[14]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _085_ (.ZN(la_data_out[15]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _086_ (.ZN(la_data_out[16]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _087_ (.ZN(la_data_out[17]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _088_ (.ZN(la_data_out[18]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _089_ (.ZN(la_data_out[19]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _090_ (.ZN(la_data_out[20]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _091_ (.ZN(la_data_out[21]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _092_ (.ZN(la_data_out[22]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _093_ (.ZN(la_data_out[23]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _094_ (.ZN(la_data_out[24]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _095_ (.ZN(la_data_out[25]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _096_ (.ZN(la_data_out[26]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _097_ (.ZN(la_data_out[27]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _098_ (.ZN(la_data_out[28]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _099_ (.ZN(la_data_out[29]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _100_ (.ZN(la_data_out[30]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _101_ (.ZN(la_data_out[31]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _102_ (.ZN(la_data_out[32]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _103_ (.ZN(la_data_out[33]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _104_ (.ZN(la_data_out[34]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _105_ (.ZN(la_data_out[35]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _106_ (.ZN(la_data_out[36]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _107_ (.ZN(la_data_out[37]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _108_ (.ZN(la_data_out[38]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _109_ (.ZN(la_data_out[39]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _110_ (.ZN(la_data_out[40]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _111_ (.ZN(la_data_out[41]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _112_ (.ZN(la_data_out[42]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _113_ (.ZN(la_data_out[43]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _114_ (.ZN(la_data_out[44]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _115_ (.ZN(la_data_out[45]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _116_ (.ZN(la_data_out[46]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _117_ (.ZN(la_data_out[47]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _118_ (.ZN(la_data_out[48]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _119_ (.ZN(la_data_out[49]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _120_ (.ZN(la_data_out[50]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _121_ (.ZN(la_data_out[51]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _122_ (.ZN(la_data_out[52]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _123_ (.ZN(la_data_out[53]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _124_ (.ZN(la_data_out[54]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _125_ (.ZN(la_data_out[55]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _126_ (.ZN(la_data_out[56]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _127_ (.ZN(la_data_out[57]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _128_ (.ZN(la_data_out[58]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _129_ (.ZN(la_data_out[59]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _130_ (.ZN(la_data_out[60]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _131_ (.ZN(la_data_out[61]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _132_ (.ZN(la_data_out[62]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _133_ (.ZN(la_data_out[63]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _134_ (.ZN(la_data_out[64]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _135_ (.ZN(la_data_out[65]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _136_ (.ZN(la_data_out[66]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _137_ (.ZN(la_data_out[67]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _138_ (.ZN(la_data_out[68]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _139_ (.ZN(la_data_out[69]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _140_ (.ZN(la_data_out[70]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _141_ (.ZN(la_data_out[71]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _142_ (.ZN(la_data_out[72]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _143_ (.ZN(la_data_out[73]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _144_ (.ZN(la_data_out[74]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _145_ (.ZN(la_data_out[75]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _146_ (.ZN(la_data_out[76]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _147_ (.ZN(la_data_out[77]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _148_ (.ZN(la_data_out[78]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _149_ (.ZN(la_data_out[79]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _150_ (.ZN(la_data_out[80]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _151_ (.ZN(la_data_out[81]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _152_ (.ZN(la_data_out[82]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _153_ (.ZN(la_data_out[83]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _154_ (.ZN(la_data_out[84]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _155_ (.ZN(la_data_out[85]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _156_ (.ZN(la_data_out[86]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _157_ (.ZN(la_data_out[87]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _158_ (.ZN(la_data_out[88]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _159_ (.ZN(la_data_out[89]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _160_ (.ZN(la_data_out[90]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _161_ (.ZN(la_data_out[91]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _162_ (.ZN(la_data_out[92]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _163_ (.ZN(la_data_out[93]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _164_ (.ZN(la_data_out[94]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _165_ (.ZN(la_data_out[95]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _166_ (.ZN(la_data_out[96]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _167_ (.ZN(la_data_out[97]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _168_ (.ZN(la_data_out[98]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _169_ (.ZN(la_data_out[99]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _170_ (.ZN(la_data_out[100]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _171_ (.ZN(la_data_out[101]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _172_ (.ZN(la_data_out[102]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _173_ (.ZN(la_data_out[103]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _174_ (.ZN(la_data_out[104]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _175_ (.ZN(la_data_out[105]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _176_ (.ZN(la_data_out[106]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _177_ (.ZN(la_data_out[107]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _178_ (.ZN(la_data_out[108]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _179_ (.ZN(la_data_out[109]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _180_ (.ZN(la_data_out[110]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _181_ (.ZN(la_data_out[111]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _182_ (.ZN(la_data_out[112]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _183_ (.ZN(la_data_out[113]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _184_ (.ZN(la_data_out[114]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _185_ (.ZN(la_data_out[115]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _186_ (.ZN(la_data_out[116]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _187_ (.ZN(la_data_out[117]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _188_ (.ZN(la_data_out[118]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _189_ (.ZN(la_data_out[119]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _190_ (.ZN(la_data_out[120]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _191_ (.ZN(la_data_out[121]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _192_ (.ZN(la_data_out[122]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _193_ (.ZN(la_data_out[123]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _194_ (.ZN(la_data_out[124]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _195_ (.ZN(la_data_out[125]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _196_ (.ZN(la_data_out[126]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _197_ (.ZN(la_data_out[127]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _198_ (.ZN(wbs_dat_o[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _199_ (.ZN(wbs_dat_o[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _200_ (.ZN(wbs_dat_o[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _201_ (.ZN(wbs_dat_o[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _202_ (.ZN(wbs_dat_o[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _203_ (.ZN(wbs_dat_o[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _204_ (.ZN(wbs_dat_o[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _205_ (.ZN(wbs_dat_o[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _206_ (.ZN(wbs_dat_o[8]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _207_ (.ZN(wbs_dat_o[9]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _208_ (.ZN(wbs_dat_o[10]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _209_ (.ZN(wbs_dat_o[11]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _210_ (.ZN(wbs_dat_o[12]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _211_ (.ZN(wbs_dat_o[13]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _212_ (.ZN(wbs_dat_o[14]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _213_ (.ZN(wbs_dat_o[15]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _214_ (.ZN(wbs_dat_o[16]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _215_ (.ZN(wbs_dat_o[17]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _216_ (.ZN(wbs_dat_o[18]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _217_ (.ZN(wbs_dat_o[19]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _218_ (.ZN(wbs_dat_o[20]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _219_ (.ZN(wbs_dat_o[21]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _220_ (.ZN(wbs_dat_o[22]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _221_ (.ZN(wbs_dat_o[23]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _222_ (.ZN(wbs_dat_o[24]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _223_ (.ZN(wbs_dat_o[25]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _224_ (.ZN(wbs_dat_o[26]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _225_ (.ZN(wbs_dat_o[27]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _226_ (.ZN(wbs_dat_o[28]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _227_ (.ZN(wbs_dat_o[29]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _228_ (.ZN(wbs_dat_o[30]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _229_ (.ZN(wbs_dat_o[31]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _230_ (.ZN(io_oeb[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _231_ (.ZN(io_oeb[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _232_ (.ZN(io_oeb[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _233_ (.ZN(io_oeb[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _234_ (.ZN(io_oeb[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _235_ (.ZN(io_oeb[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _236_ (.ZN(io_oeb[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _237_ (.ZN(io_oeb[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _238_ (.ZN(io_oeb[8]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__tiel _239_ (.ZN(io_oeb[9]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Right_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Right_49 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Right_50 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Right_51 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Right_52 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Right_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Right_54 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Right_55 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Right_56 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Right_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Right_58 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Right_59 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Right_60 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Right_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Right_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Right_63 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Right_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Right_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Right_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Right_67 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Right_68 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Right_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Right_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Right_71 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Right_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Right_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Right_74 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Right_75 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Right_76 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Right_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Right_78 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Right_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Right_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Right_81 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Right_82 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Right_83 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Right_84 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Right_85 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Right_86 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Right_87 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Right_88 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Right_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Right_90 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Right_91 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Right_92 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Right_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Right_94 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Right_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Right_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Right_97 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Right_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Right_99 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Right_100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Right_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Right_102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Right_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Right_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Right_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Right_106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Right_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Right_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Right_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Right_110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Right_111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Right_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Right_113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Right_114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Right_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Right_116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Right_117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Right_118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Right_119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Right_120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Right_121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Right_122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Right_123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Right_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Right_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Right_126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Right_127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Right_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Right_129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Right_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Right_131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Right_132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Right_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Right_134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Right_135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Right_136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Right_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Right_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Right_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Right_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Right_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Right_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Right_143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Right_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Right_145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Right_146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Right_147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Right_148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Right_149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Right_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Right_151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Right_152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Right_153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Right_154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Right_155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Right_156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Right_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Right_158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Right_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Right_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Right_161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Right_162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_163_Right_163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_164_Right_164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_165_Right_165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_166_Right_166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_167_Right_167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_168_Right_168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_169_Right_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_170_Right_170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_171_Right_171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_172_Right_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_173_Right_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_174_Right_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_175_Right_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_176_Right_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_177_Right_177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_178_Right_178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_179_Right_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_180_Right_180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_181_Right_181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_182_Right_182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_183_Right_183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_184_Right_184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_185_Right_185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_186_Right_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_187_Right_187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_188_Right_188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_189_Right_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_190_Right_190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_191_Right_191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_192_Right_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_193_Right_193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_194_Right_194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_195_Right_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_196_Right_196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_197_Right_197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_198_Right_198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_199_Right_199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_200_Right_200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_201_Right_201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_202_Right_202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_203_Right_203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_204_Right_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_205_Right_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_206_Right_206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_207_Right_207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_208_Right_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_209_Right_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_210_Right_210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_211_Right_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_212_Right_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_213_Right_213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_214_Right_214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_215_Right_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_216_Right_216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_217_Right_217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_218_Right_218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_219_Right_219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_220_Right_220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_221_Right_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_222_Right_222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_223_Right_223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_224_Right_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_225_Right_225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_226_Right_226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_227_Right_227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_228_Right_228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_229_Right_229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_230_Right_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_231_Right_231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_232_Right_232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_233_Right_233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_234_Right_234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_235_Right_235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_236_Right_236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_237_Right_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_238_Right_238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_239_Right_239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_240_Right_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_241_Right_241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_242_Right_242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_243_Right_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_244_Right_244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_245_Right_245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_246_Right_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_247_Right_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_248_Right_248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_249_Right_249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_250_Right_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_251_Right_251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_252_Right_252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_253_Right_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_254_Right_254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_255_Right_255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_256_Right_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_257_Right_257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_258_Right_258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_259_Right_259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_260_Right_260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_261_Right_261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_262_Right_262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_263_Right_263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_264_Right_264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_265_Right_265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_266_Right_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_267_Right_267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_268_Right_268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_269_Right_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_270_Right_270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_271_Right_271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_272_Right_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_273_Right_273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_274_Right_274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_275_Right_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_276_Right_276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_277_Right_277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_278_Right_278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_279_Right_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_280_Right_280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_281_Right_281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_282_Right_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_283_Right_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_284_Right_284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_285_Right_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_286_Right_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_287_Right_287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_288_Right_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_289_Right_289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_290_Right_290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_291_Right_291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_292_Right_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_293_Right_293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_294_Right_294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_295_Right_295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_296_Right_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_297_Right_297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_298_Right_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_299_Right_299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_300_Right_300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_301_Right_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_302_Right_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_303_Right_303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_304_Right_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_305_Right_305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_306_Right_306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_307_Right_307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_308_Right_308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_309_Right_309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_310_Right_310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_311_Right_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_312_Right_312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_313_Right_313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_314_Right_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_315_Right_315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_316_Right_316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_317_Right_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_318_Right_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_319_Right_319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_320_Right_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_321_Right_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_322_Right_322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_323_Right_323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_324_Right_324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_325_Right_325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_326_Right_326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_327_Right_327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_328_Right_328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_329_Right_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_330_Right_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_331_Right_331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_332_Right_332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_333_Right_333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_334_Right_334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_335_Right_335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_336_Right_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_337_Right_337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_338_Right_338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_339_Right_339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_340_Right_340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_341_Right_341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Left_390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Left_391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Left_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Left_393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Left_394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Left_395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Left_396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Left_397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Left_398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Left_399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Left_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Left_401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Left_402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Left_403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Left_404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Left_405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Left_406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Left_407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Left_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Left_409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Left_410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Left_411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Left_412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Left_413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Left_414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Left_415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Left_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Left_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Left_418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Left_419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Left_420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Left_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Left_422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Left_423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Left_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Left_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Left_426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Left_427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Left_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Left_429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Left_430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Left_431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Left_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Left_433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Left_434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Left_435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Left_436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Left_437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Left_438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Left_439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Left_440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Left_441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Left_442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Left_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Left_444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_103_Left_445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_104_Left_446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_105_Left_447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_106_Left_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_107_Left_449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_108_Left_450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_109_Left_451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_110_Left_452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_111_Left_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_112_Left_454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_113_Left_455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_114_Left_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_115_Left_457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_116_Left_458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_117_Left_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_118_Left_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_119_Left_461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_120_Left_462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_121_Left_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_122_Left_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_123_Left_465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_124_Left_466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_125_Left_467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_126_Left_468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_127_Left_469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_128_Left_470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_129_Left_471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_130_Left_472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_131_Left_473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_132_Left_474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_133_Left_475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_134_Left_476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_135_Left_477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_136_Left_478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_137_Left_479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_138_Left_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_139_Left_481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_140_Left_482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_141_Left_483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_142_Left_484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_143_Left_485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_144_Left_486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_145_Left_487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_146_Left_488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_147_Left_489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_148_Left_490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_149_Left_491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_150_Left_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_151_Left_493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_152_Left_494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_153_Left_495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_154_Left_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_155_Left_497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_156_Left_498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_157_Left_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_158_Left_500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_159_Left_501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_160_Left_502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_161_Left_503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_162_Left_504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_163_Left_505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_164_Left_506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_165_Left_507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_166_Left_508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_167_Left_509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_168_Left_510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_169_Left_511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_170_Left_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_171_Left_513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_172_Left_514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_173_Left_515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_174_Left_516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_175_Left_517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_176_Left_518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_177_Left_519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_178_Left_520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_179_Left_521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_180_Left_522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_181_Left_523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_182_Left_524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_183_Left_525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_184_Left_526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_185_Left_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_186_Left_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_187_Left_529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_188_Left_530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_189_Left_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_190_Left_532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_191_Left_533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_192_Left_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_193_Left_535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_194_Left_536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_195_Left_537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_196_Left_538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_197_Left_539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_198_Left_540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_199_Left_541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_200_Left_542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_201_Left_543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_202_Left_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_203_Left_545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_204_Left_546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_205_Left_547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_206_Left_548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_207_Left_549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_208_Left_550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_209_Left_551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_210_Left_552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_211_Left_553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_212_Left_554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_213_Left_555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_214_Left_556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_215_Left_557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_216_Left_558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_217_Left_559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_218_Left_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_219_Left_561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_220_Left_562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_221_Left_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_222_Left_564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_223_Left_565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_224_Left_566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_225_Left_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_226_Left_568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_227_Left_569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_228_Left_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_229_Left_571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_230_Left_572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_231_Left_573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_232_Left_574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_233_Left_575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_234_Left_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_235_Left_577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_236_Left_578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_237_Left_579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_238_Left_580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_239_Left_581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_240_Left_582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_241_Left_583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_242_Left_584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_243_Left_585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_244_Left_586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_245_Left_587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_246_Left_588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_247_Left_589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_248_Left_590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_249_Left_591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_250_Left_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_251_Left_593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_252_Left_594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_253_Left_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_254_Left_596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_255_Left_597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_256_Left_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_257_Left_599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_258_Left_600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_259_Left_601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_260_Left_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_261_Left_603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_262_Left_604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_263_Left_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_264_Left_606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_265_Left_607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_266_Left_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_267_Left_609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_268_Left_610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_269_Left_611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_270_Left_612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_271_Left_613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_272_Left_614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_273_Left_615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_274_Left_616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_275_Left_617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_276_Left_618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_277_Left_619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_278_Left_620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_279_Left_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_280_Left_622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_281_Left_623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_282_Left_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_283_Left_625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_284_Left_626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_285_Left_627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_286_Left_628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_287_Left_629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_288_Left_630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_289_Left_631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_290_Left_632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_291_Left_633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_292_Left_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_293_Left_635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_294_Left_636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_295_Left_637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_296_Left_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_297_Left_639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_298_Left_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_299_Left_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_300_Left_642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_301_Left_643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_302_Left_644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_303_Left_645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_304_Left_646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_305_Left_647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_306_Left_648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_307_Left_649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_308_Left_650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_309_Left_651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_310_Left_652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_311_Left_653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_312_Left_654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_313_Left_655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_314_Left_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_315_Left_657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_316_Left_658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_317_Left_659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_318_Left_660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_319_Left_661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_320_Left_662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_321_Left_663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_322_Left_664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_323_Left_665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_324_Left_666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_325_Left_667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_326_Left_668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_327_Left_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_328_Left_670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_329_Left_671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_330_Left_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_331_Left_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_332_Left_674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_333_Left_675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_334_Left_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_335_Left_677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_336_Left_678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_337_Left_679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_338_Left_680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_339_Left_681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_340_Left_682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_341_Left_683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_1042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_1113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_1255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_1326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_1397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_1468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_1539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_1610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_1681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_1752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_1823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_1894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_1965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_1999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_2036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_2107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_2178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_2249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_2391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_2462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_2533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_2604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_2675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_2746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_2817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_2888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_2959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_2999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_3030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_3101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_3172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_3243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_3314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_3385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_3527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_3598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_3669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_3740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_3811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_3882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_3953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_3999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_4024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_4095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_4166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_4237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_4308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_4379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_4450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_4521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_4663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_4734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_4805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_4876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_4947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_4999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_5000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_5001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_5002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_5003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_5004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_5005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_5006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_5007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_5009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_5010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_5011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_5012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_5013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_5014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_5015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_5016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_5017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_5018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_5089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_5160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_5231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_5302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_5373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_5444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_5515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_5586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_5657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_5799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_5870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_5941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_5999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_6001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_6002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_6003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_6004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_6005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_6006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_6007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_6008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_6009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_6010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_6011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_6012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_6083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_6154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_6225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_6296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_6367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_6438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_6509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_6580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_6651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_6722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_6793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_6935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_6999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_7000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_7001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_7002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_7003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_7004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_7005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_7006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_7077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_7148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_7219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_7290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_7361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_7432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_7503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_7574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_7645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_7716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_7787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_7858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_7929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_7999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_8071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_103_8142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_104_8213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_105_8284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_106_8355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_107_8426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_108_8497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_109_8568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_110_8639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_111_8710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_112_8781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_113_8852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_114_8923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_115_8994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_8995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_8996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_8997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_8998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_8999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_116_9065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_117_9136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_118_9207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_119_9278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_120_9349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_121_9420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_122_9491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_123_9562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_124_9633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_125_9704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_126_9775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_127_9846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_128_9917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_129_9988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_9989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_9990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_9991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_9992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_9993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_9994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_9995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_9996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_9997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_9998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_9999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_130_10059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_131_10130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_132_10201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_133_10272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_134_10343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_135_10414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_136_10485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_137_10556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_138_10627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_139_10698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_140_10769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_141_10840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_142_10911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_143_10982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_10983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_10984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_10985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_10986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_10987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_10988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_10989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_10990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_10991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_10992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_10993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_10994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_10995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_10996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_10997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_10998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_10999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_144_11053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_145_11124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_146_11195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_147_11266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_148_11337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_149_11408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_150_11479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_151_11550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_152_11621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_153_11692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_154_11763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_155_11834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_156_11905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_157_11976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_11999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_158_12047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_159_12118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_160_12189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_161_12260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_162_12331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_163_12402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_164_12473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_165_12544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_166_12615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_167_12686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_168_12757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_169_12828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_170_12899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_171_12970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_12999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_172_13041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_173_13112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_174_13183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_175_13254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_176_13325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_177_13396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_178_13467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_179_13538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_180_13609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_181_13680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_182_13751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_183_13822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_184_13893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_185_13964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_13999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_186_14035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_187_14106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_188_14177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_189_14248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_190_14319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_191_14390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_192_14461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_193_14532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_194_14603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_195_14674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_196_14745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_197_14816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_198_14887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_199_14958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_14999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_200_15029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_201_15100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_202_15171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_203_15242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_204_15313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_205_15384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_206_15455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_207_15526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_208_15597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_209_15668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_210_15739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_211_15810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_212_15881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_213_15952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_15999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_214_16023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_215_16094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_216_16165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_217_16236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_218_16307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_219_16378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_220_16449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_221_16520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_222_16591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_223_16662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_224_16733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_225_16804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_226_16875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_227_16946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_16999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_17000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_17001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_17002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_17003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_17004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_17005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_17006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_17007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_17008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_17009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_17010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_17011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_17012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_17013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_17014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_17015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_17016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_228_17017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_229_17088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_230_17159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_231_17230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_232_17301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_233_17372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_234_17443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_235_17514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_236_17585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_237_17656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_238_17727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_239_17798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_240_17869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_241_17940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_17999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_18000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_18001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_18002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_18003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_18004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_18005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_18006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_18007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_18008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_18009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_18010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_242_18011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_243_18082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_244_18153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_245_18224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_246_18295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_247_18366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_248_18437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_249_18508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_250_18579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_251_18650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_252_18721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_253_18792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_254_18863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_255_18934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_18999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_19000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_19001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_19002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_19003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_19004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_256_19005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_257_19076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_258_19147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_259_19218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_260_19289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_261_19360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_262_19431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_263_19502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_264_19573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_265_19644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_266_19715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_267_19786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_268_19857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_269_19928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_270_19999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_271_20070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_272_20141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_273_20212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_274_20283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_275_20354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_276_20425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_277_20496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_278_20567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_279_20638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_280_20709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_281_20780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_282_20851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_283_20922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_284_20993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_20994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_20995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_20996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_20997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_20998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_20999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_285_21064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_286_21135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_287_21206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_288_21277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_289_21348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_290_21419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_291_21490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_292_21561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_293_21632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_294_21703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_295_21774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_296_21845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_297_21916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_298_21987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_21988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_21989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_21990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_21991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_21992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_21993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_21994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_21995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_21996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_21997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_21998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_21999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_299_22058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_300_22129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_301_22200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_302_22271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_303_22342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_304_22413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_305_22484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_306_22555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_307_22626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_308_22697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_309_22768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_310_22839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_311_22910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_312_22981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_22982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_22983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_22984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_22985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_22986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_22987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_22988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_22989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_22990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_22991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_22992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_22993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_22994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_22995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_22996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_22997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_22998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_22999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_313_23052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_314_23123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_315_23194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_316_23265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_317_23336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_318_23407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_319_23478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_320_23549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_321_23620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_322_23691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_323_23762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_324_23833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_325_23904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_326_23975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_23999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_327_24046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_328_24117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_329_24188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_330_24259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_331_24330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_332_24401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_333_24472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_334_24543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_335_24614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_336_24685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_337_24756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_338_24827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_339_24898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_340_24969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_24999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_341_25115 (.VDD(vdd),
    .VSS(vss));
endmodule
